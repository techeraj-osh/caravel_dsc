magic
tech sky130A
magscale 1 2
timestamp 1623609253
<< obsli1 >>
rect 1104 2159 111136 112081
<< obsm1 >>
rect 106 1028 112226 112112
<< metal2 >>
rect 478 113654 534 114454
rect 1398 113654 1454 114454
rect 2410 113654 2466 114454
rect 3422 113654 3478 114454
rect 4342 113654 4398 114454
rect 5354 113654 5410 114454
rect 6366 113654 6422 114454
rect 7286 113654 7342 114454
rect 8298 113654 8354 114454
rect 9310 113654 9366 114454
rect 10322 113654 10378 114454
rect 11242 113654 11298 114454
rect 12254 113654 12310 114454
rect 13266 113654 13322 114454
rect 14186 113654 14242 114454
rect 15198 113654 15254 114454
rect 16210 113654 16266 114454
rect 17222 113654 17278 114454
rect 18142 113654 18198 114454
rect 19154 113654 19210 114454
rect 20166 113654 20222 114454
rect 21086 113654 21142 114454
rect 22098 113654 22154 114454
rect 23110 113654 23166 114454
rect 24122 113654 24178 114454
rect 25042 113654 25098 114454
rect 26054 113654 26110 114454
rect 27066 113654 27122 114454
rect 27986 113654 28042 114454
rect 28998 113654 29054 114454
rect 30010 113654 30066 114454
rect 31022 113654 31078 114454
rect 31942 113654 31998 114454
rect 32954 113654 33010 114454
rect 33966 113654 34022 114454
rect 34886 113654 34942 114454
rect 35898 113654 35954 114454
rect 36910 113654 36966 114454
rect 37922 113654 37978 114454
rect 38842 113654 38898 114454
rect 39854 113654 39910 114454
rect 40866 113654 40922 114454
rect 41786 113654 41842 114454
rect 42798 113654 42854 114454
rect 43810 113654 43866 114454
rect 44730 113654 44786 114454
rect 45742 113654 45798 114454
rect 46754 113654 46810 114454
rect 47766 113654 47822 114454
rect 48686 113654 48742 114454
rect 49698 113654 49754 114454
rect 50710 113654 50766 114454
rect 51630 113654 51686 114454
rect 52642 113654 52698 114454
rect 53654 113654 53710 114454
rect 54666 113654 54722 114454
rect 55586 113654 55642 114454
rect 56598 113654 56654 114454
rect 57610 113654 57666 114454
rect 58530 113654 58586 114454
rect 59542 113654 59598 114454
rect 60554 113654 60610 114454
rect 61566 113654 61622 114454
rect 62486 113654 62542 114454
rect 63498 113654 63554 114454
rect 64510 113654 64566 114454
rect 65430 113654 65486 114454
rect 66442 113654 66498 114454
rect 67454 113654 67510 114454
rect 68466 113654 68522 114454
rect 69386 113654 69442 114454
rect 70398 113654 70454 114454
rect 71410 113654 71466 114454
rect 72330 113654 72386 114454
rect 73342 113654 73398 114454
rect 74354 113654 74410 114454
rect 75366 113654 75422 114454
rect 76286 113654 76342 114454
rect 77298 113654 77354 114454
rect 78310 113654 78366 114454
rect 79230 113654 79286 114454
rect 80242 113654 80298 114454
rect 81254 113654 81310 114454
rect 82174 113654 82230 114454
rect 83186 113654 83242 114454
rect 84198 113654 84254 114454
rect 85210 113654 85266 114454
rect 86130 113654 86186 114454
rect 87142 113654 87198 114454
rect 88154 113654 88210 114454
rect 89074 113654 89130 114454
rect 90086 113654 90142 114454
rect 91098 113654 91154 114454
rect 92110 113654 92166 114454
rect 93030 113654 93086 114454
rect 94042 113654 94098 114454
rect 95054 113654 95110 114454
rect 95974 113654 96030 114454
rect 96986 113654 97042 114454
rect 97998 113654 98054 114454
rect 99010 113654 99066 114454
rect 99930 113654 99986 114454
rect 100942 113654 100998 114454
rect 101954 113654 102010 114454
rect 102874 113654 102930 114454
rect 103886 113654 103942 114454
rect 104898 113654 104954 114454
rect 105910 113654 105966 114454
rect 106830 113654 106886 114454
rect 107842 113654 107898 114454
rect 108854 113654 108910 114454
rect 109774 113654 109830 114454
rect 110786 113654 110842 114454
rect 111798 113654 111854 114454
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 754 0 810 800
rect 938 0 994 800
rect 1214 0 1270 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2318 0 2374 800
rect 2594 0 2650 800
rect 2778 0 2834 800
rect 3054 0 3110 800
rect 3238 0 3294 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5814 0 5870 800
rect 5998 0 6054 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7654 0 7710 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8758 0 8814 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10138 0 10194 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11334 0 11390 800
rect 11518 0 11574 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 13174 0 13230 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 14922 0 14978 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15658 0 15714 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16578 0 16634 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19338 0 19394 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20442 0 20498 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22282 0 22338 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 25962 0 26018 800
rect 26238 0 26294 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27618 0 27674 800
rect 27802 0 27858 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28446 0 28502 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29826 0 29882 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31206 0 31262 800
rect 31482 0 31538 800
rect 31666 0 31722 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32862 0 32918 800
rect 33046 0 33102 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 37002 0 37058 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38842 0 38898 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39762 0 39818 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41602 0 41658 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44730 0 44786 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48226 0 48282 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49606 0 49662 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51630 0 51686 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52366 0 52422 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53746 0 53802 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56690 0 56746 800
rect 56874 0 56930 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58530 0 58586 800
rect 58714 0 58770 800
rect 58990 0 59046 800
rect 59174 0 59230 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59910 0 59966 800
rect 60094 0 60150 800
rect 60370 0 60426 800
rect 60554 0 60610 800
rect 60830 0 60886 800
rect 61014 0 61070 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62210 0 62266 800
rect 62394 0 62450 800
rect 62670 0 62726 800
rect 62854 0 62910 800
rect 63130 0 63186 800
rect 63314 0 63370 800
rect 63590 0 63646 800
rect 63774 0 63830 800
rect 64050 0 64106 800
rect 64234 0 64290 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64970 0 65026 800
rect 65154 0 65210 800
rect 65430 0 65486 800
rect 65614 0 65670 800
rect 65890 0 65946 800
rect 66074 0 66130 800
rect 66350 0 66406 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 66994 0 67050 800
rect 67270 0 67326 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68650 0 68706 800
rect 68834 0 68890 800
rect 69110 0 69166 800
rect 69294 0 69350 800
rect 69570 0 69626 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70214 0 70270 800
rect 70398 0 70454 800
rect 70674 0 70730 800
rect 70858 0 70914 800
rect 71134 0 71190 800
rect 71318 0 71374 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72514 0 72570 800
rect 72698 0 72754 800
rect 72974 0 73030 800
rect 73158 0 73214 800
rect 73434 0 73490 800
rect 73618 0 73674 800
rect 73894 0 73950 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74538 0 74594 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76378 0 76434 800
rect 76654 0 76710 800
rect 76838 0 76894 800
rect 77114 0 77170 800
rect 77298 0 77354 800
rect 77574 0 77630 800
rect 77758 0 77814 800
rect 78034 0 78090 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78954 0 79010 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79598 0 79654 800
rect 79874 0 79930 800
rect 80058 0 80114 800
rect 80334 0 80390 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 80978 0 81034 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 81898 0 81954 800
rect 82174 0 82230 800
rect 82358 0 82414 800
rect 82634 0 82690 800
rect 82818 0 82874 800
rect 83094 0 83150 800
rect 83278 0 83334 800
rect 83554 0 83610 800
rect 83738 0 83794 800
rect 84014 0 84070 800
rect 84198 0 84254 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84842 0 84898 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85578 0 85634 800
rect 85762 0 85818 800
rect 86038 0 86094 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86682 0 86738 800
rect 86958 0 87014 800
rect 87142 0 87198 800
rect 87418 0 87474 800
rect 87602 0 87658 800
rect 87878 0 87934 800
rect 88062 0 88118 800
rect 88338 0 88394 800
rect 88522 0 88578 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89258 0 89314 800
rect 89442 0 89498 800
rect 89718 0 89774 800
rect 89902 0 89958 800
rect 90178 0 90234 800
rect 90362 0 90418 800
rect 90638 0 90694 800
rect 90822 0 90878 800
rect 91098 0 91154 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 92018 0 92074 800
rect 92202 0 92258 800
rect 92478 0 92534 800
rect 92662 0 92718 800
rect 92938 0 92994 800
rect 93122 0 93178 800
rect 93398 0 93454 800
rect 93582 0 93638 800
rect 93858 0 93914 800
rect 94042 0 94098 800
rect 94318 0 94374 800
rect 94502 0 94558 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95698 0 95754 800
rect 95882 0 95938 800
rect 96158 0 96214 800
rect 96342 0 96398 800
rect 96618 0 96674 800
rect 96802 0 96858 800
rect 97078 0 97134 800
rect 97262 0 97318 800
rect 97538 0 97594 800
rect 97722 0 97778 800
rect 97998 0 98054 800
rect 98182 0 98238 800
rect 98366 0 98422 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99102 0 99158 800
rect 99286 0 99342 800
rect 99562 0 99618 800
rect 99746 0 99802 800
rect 100022 0 100078 800
rect 100206 0 100262 800
rect 100482 0 100538 800
rect 100666 0 100722 800
rect 100942 0 100998 800
rect 101126 0 101182 800
rect 101402 0 101458 800
rect 101586 0 101642 800
rect 101862 0 101918 800
rect 102046 0 102102 800
rect 102322 0 102378 800
rect 102506 0 102562 800
rect 102782 0 102838 800
rect 102966 0 103022 800
rect 103242 0 103298 800
rect 103426 0 103482 800
rect 103702 0 103758 800
rect 103886 0 103942 800
rect 104162 0 104218 800
rect 104346 0 104402 800
rect 104622 0 104678 800
rect 104806 0 104862 800
rect 105082 0 105138 800
rect 105266 0 105322 800
rect 105542 0 105598 800
rect 105726 0 105782 800
rect 106002 0 106058 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106646 0 106702 800
rect 106922 0 106978 800
rect 107106 0 107162 800
rect 107382 0 107438 800
rect 107566 0 107622 800
rect 107842 0 107898 800
rect 108026 0 108082 800
rect 108302 0 108358 800
rect 108486 0 108542 800
rect 108762 0 108818 800
rect 108946 0 109002 800
rect 109222 0 109278 800
rect 109406 0 109462 800
rect 109682 0 109738 800
rect 109866 0 109922 800
rect 110142 0 110198 800
rect 110326 0 110382 800
rect 110602 0 110658 800
rect 110786 0 110842 800
rect 111062 0 111118 800
rect 111246 0 111302 800
rect 111522 0 111578 800
rect 111706 0 111762 800
rect 111982 0 112038 800
rect 112166 0 112222 800
<< obsm2 >>
rect 112 113598 422 113654
rect 590 113598 1342 113654
rect 1510 113598 2354 113654
rect 2522 113598 3366 113654
rect 3534 113598 4286 113654
rect 4454 113598 5298 113654
rect 5466 113598 6310 113654
rect 6478 113598 7230 113654
rect 7398 113598 8242 113654
rect 8410 113598 9254 113654
rect 9422 113598 10266 113654
rect 10434 113598 11186 113654
rect 11354 113598 12198 113654
rect 12366 113598 13210 113654
rect 13378 113598 14130 113654
rect 14298 113598 15142 113654
rect 15310 113598 16154 113654
rect 16322 113598 17166 113654
rect 17334 113598 18086 113654
rect 18254 113598 19098 113654
rect 19266 113598 20110 113654
rect 20278 113598 21030 113654
rect 21198 113598 22042 113654
rect 22210 113598 23054 113654
rect 23222 113598 24066 113654
rect 24234 113598 24986 113654
rect 25154 113598 25998 113654
rect 26166 113598 27010 113654
rect 27178 113598 27930 113654
rect 28098 113598 28942 113654
rect 29110 113598 29954 113654
rect 30122 113598 30966 113654
rect 31134 113598 31886 113654
rect 32054 113598 32898 113654
rect 33066 113598 33910 113654
rect 34078 113598 34830 113654
rect 34998 113598 35842 113654
rect 36010 113598 36854 113654
rect 37022 113598 37866 113654
rect 38034 113598 38786 113654
rect 38954 113598 39798 113654
rect 39966 113598 40810 113654
rect 40978 113598 41730 113654
rect 41898 113598 42742 113654
rect 42910 113598 43754 113654
rect 43922 113598 44674 113654
rect 44842 113598 45686 113654
rect 45854 113598 46698 113654
rect 46866 113598 47710 113654
rect 47878 113598 48630 113654
rect 48798 113598 49642 113654
rect 49810 113598 50654 113654
rect 50822 113598 51574 113654
rect 51742 113598 52586 113654
rect 52754 113598 53598 113654
rect 53766 113598 54610 113654
rect 54778 113598 55530 113654
rect 55698 113598 56542 113654
rect 56710 113598 57554 113654
rect 57722 113598 58474 113654
rect 58642 113598 59486 113654
rect 59654 113598 60498 113654
rect 60666 113598 61510 113654
rect 61678 113598 62430 113654
rect 62598 113598 63442 113654
rect 63610 113598 64454 113654
rect 64622 113598 65374 113654
rect 65542 113598 66386 113654
rect 66554 113598 67398 113654
rect 67566 113598 68410 113654
rect 68578 113598 69330 113654
rect 69498 113598 70342 113654
rect 70510 113598 71354 113654
rect 71522 113598 72274 113654
rect 72442 113598 73286 113654
rect 73454 113598 74298 113654
rect 74466 113598 75310 113654
rect 75478 113598 76230 113654
rect 76398 113598 77242 113654
rect 77410 113598 78254 113654
rect 78422 113598 79174 113654
rect 79342 113598 80186 113654
rect 80354 113598 81198 113654
rect 81366 113598 82118 113654
rect 82286 113598 83130 113654
rect 83298 113598 84142 113654
rect 84310 113598 85154 113654
rect 85322 113598 86074 113654
rect 86242 113598 87086 113654
rect 87254 113598 88098 113654
rect 88266 113598 89018 113654
rect 89186 113598 90030 113654
rect 90198 113598 91042 113654
rect 91210 113598 92054 113654
rect 92222 113598 92974 113654
rect 93142 113598 93986 113654
rect 94154 113598 94998 113654
rect 95166 113598 95918 113654
rect 96086 113598 96930 113654
rect 97098 113598 97942 113654
rect 98110 113598 98954 113654
rect 99122 113598 99874 113654
rect 100042 113598 100886 113654
rect 101054 113598 101898 113654
rect 102066 113598 102818 113654
rect 102986 113598 103830 113654
rect 103998 113598 104842 113654
rect 105010 113598 105854 113654
rect 106022 113598 106774 113654
rect 106942 113598 107786 113654
rect 107954 113598 108798 113654
rect 108966 113598 109718 113654
rect 109886 113598 110730 113654
rect 110898 113598 111742 113654
rect 111910 113598 112220 113654
rect 112 856 112220 113598
rect 222 800 238 856
rect 406 800 422 856
rect 590 800 698 856
rect 866 800 882 856
rect 1050 800 1158 856
rect 1326 800 1342 856
rect 1510 800 1618 856
rect 1786 800 1802 856
rect 1970 800 2078 856
rect 2246 800 2262 856
rect 2430 800 2538 856
rect 2706 800 2722 856
rect 2890 800 2998 856
rect 3166 800 3182 856
rect 3350 800 3458 856
rect 3626 800 3642 856
rect 3810 800 3918 856
rect 4086 800 4102 856
rect 4270 800 4378 856
rect 4546 800 4562 856
rect 4730 800 4838 856
rect 5006 800 5022 856
rect 5190 800 5298 856
rect 5466 800 5482 856
rect 5650 800 5758 856
rect 5926 800 5942 856
rect 6110 800 6218 856
rect 6386 800 6402 856
rect 6570 800 6678 856
rect 6846 800 6862 856
rect 7030 800 7138 856
rect 7306 800 7322 856
rect 7490 800 7598 856
rect 7766 800 7782 856
rect 7950 800 8058 856
rect 8226 800 8242 856
rect 8410 800 8518 856
rect 8686 800 8702 856
rect 8870 800 8978 856
rect 9146 800 9162 856
rect 9330 800 9438 856
rect 9606 800 9622 856
rect 9790 800 9898 856
rect 10066 800 10082 856
rect 10250 800 10358 856
rect 10526 800 10542 856
rect 10710 800 10818 856
rect 10986 800 11002 856
rect 11170 800 11278 856
rect 11446 800 11462 856
rect 11630 800 11738 856
rect 11906 800 11922 856
rect 12090 800 12198 856
rect 12366 800 12382 856
rect 12550 800 12658 856
rect 12826 800 12842 856
rect 13010 800 13118 856
rect 13286 800 13302 856
rect 13470 800 13578 856
rect 13746 800 13762 856
rect 13930 800 14038 856
rect 14206 800 14222 856
rect 14390 800 14406 856
rect 14574 800 14682 856
rect 14850 800 14866 856
rect 15034 800 15142 856
rect 15310 800 15326 856
rect 15494 800 15602 856
rect 15770 800 15786 856
rect 15954 800 16062 856
rect 16230 800 16246 856
rect 16414 800 16522 856
rect 16690 800 16706 856
rect 16874 800 16982 856
rect 17150 800 17166 856
rect 17334 800 17442 856
rect 17610 800 17626 856
rect 17794 800 17902 856
rect 18070 800 18086 856
rect 18254 800 18362 856
rect 18530 800 18546 856
rect 18714 800 18822 856
rect 18990 800 19006 856
rect 19174 800 19282 856
rect 19450 800 19466 856
rect 19634 800 19742 856
rect 19910 800 19926 856
rect 20094 800 20202 856
rect 20370 800 20386 856
rect 20554 800 20662 856
rect 20830 800 20846 856
rect 21014 800 21122 856
rect 21290 800 21306 856
rect 21474 800 21582 856
rect 21750 800 21766 856
rect 21934 800 22042 856
rect 22210 800 22226 856
rect 22394 800 22502 856
rect 22670 800 22686 856
rect 22854 800 22962 856
rect 23130 800 23146 856
rect 23314 800 23422 856
rect 23590 800 23606 856
rect 23774 800 23882 856
rect 24050 800 24066 856
rect 24234 800 24342 856
rect 24510 800 24526 856
rect 24694 800 24802 856
rect 24970 800 24986 856
rect 25154 800 25262 856
rect 25430 800 25446 856
rect 25614 800 25722 856
rect 25890 800 25906 856
rect 26074 800 26182 856
rect 26350 800 26366 856
rect 26534 800 26642 856
rect 26810 800 26826 856
rect 26994 800 27102 856
rect 27270 800 27286 856
rect 27454 800 27562 856
rect 27730 800 27746 856
rect 27914 800 28022 856
rect 28190 800 28206 856
rect 28374 800 28390 856
rect 28558 800 28666 856
rect 28834 800 28850 856
rect 29018 800 29126 856
rect 29294 800 29310 856
rect 29478 800 29586 856
rect 29754 800 29770 856
rect 29938 800 30046 856
rect 30214 800 30230 856
rect 30398 800 30506 856
rect 30674 800 30690 856
rect 30858 800 30966 856
rect 31134 800 31150 856
rect 31318 800 31426 856
rect 31594 800 31610 856
rect 31778 800 31886 856
rect 32054 800 32070 856
rect 32238 800 32346 856
rect 32514 800 32530 856
rect 32698 800 32806 856
rect 32974 800 32990 856
rect 33158 800 33266 856
rect 33434 800 33450 856
rect 33618 800 33726 856
rect 33894 800 33910 856
rect 34078 800 34186 856
rect 34354 800 34370 856
rect 34538 800 34646 856
rect 34814 800 34830 856
rect 34998 800 35106 856
rect 35274 800 35290 856
rect 35458 800 35566 856
rect 35734 800 35750 856
rect 35918 800 36026 856
rect 36194 800 36210 856
rect 36378 800 36486 856
rect 36654 800 36670 856
rect 36838 800 36946 856
rect 37114 800 37130 856
rect 37298 800 37406 856
rect 37574 800 37590 856
rect 37758 800 37866 856
rect 38034 800 38050 856
rect 38218 800 38326 856
rect 38494 800 38510 856
rect 38678 800 38786 856
rect 38954 800 38970 856
rect 39138 800 39246 856
rect 39414 800 39430 856
rect 39598 800 39706 856
rect 39874 800 39890 856
rect 40058 800 40166 856
rect 40334 800 40350 856
rect 40518 800 40626 856
rect 40794 800 40810 856
rect 40978 800 41086 856
rect 41254 800 41270 856
rect 41438 800 41546 856
rect 41714 800 41730 856
rect 41898 800 42006 856
rect 42174 800 42190 856
rect 42358 800 42374 856
rect 42542 800 42650 856
rect 42818 800 42834 856
rect 43002 800 43110 856
rect 43278 800 43294 856
rect 43462 800 43570 856
rect 43738 800 43754 856
rect 43922 800 44030 856
rect 44198 800 44214 856
rect 44382 800 44490 856
rect 44658 800 44674 856
rect 44842 800 44950 856
rect 45118 800 45134 856
rect 45302 800 45410 856
rect 45578 800 45594 856
rect 45762 800 45870 856
rect 46038 800 46054 856
rect 46222 800 46330 856
rect 46498 800 46514 856
rect 46682 800 46790 856
rect 46958 800 46974 856
rect 47142 800 47250 856
rect 47418 800 47434 856
rect 47602 800 47710 856
rect 47878 800 47894 856
rect 48062 800 48170 856
rect 48338 800 48354 856
rect 48522 800 48630 856
rect 48798 800 48814 856
rect 48982 800 49090 856
rect 49258 800 49274 856
rect 49442 800 49550 856
rect 49718 800 49734 856
rect 49902 800 50010 856
rect 50178 800 50194 856
rect 50362 800 50470 856
rect 50638 800 50654 856
rect 50822 800 50930 856
rect 51098 800 51114 856
rect 51282 800 51390 856
rect 51558 800 51574 856
rect 51742 800 51850 856
rect 52018 800 52034 856
rect 52202 800 52310 856
rect 52478 800 52494 856
rect 52662 800 52770 856
rect 52938 800 52954 856
rect 53122 800 53230 856
rect 53398 800 53414 856
rect 53582 800 53690 856
rect 53858 800 53874 856
rect 54042 800 54150 856
rect 54318 800 54334 856
rect 54502 800 54610 856
rect 54778 800 54794 856
rect 54962 800 55070 856
rect 55238 800 55254 856
rect 55422 800 55530 856
rect 55698 800 55714 856
rect 55882 800 55990 856
rect 56158 800 56174 856
rect 56342 800 56358 856
rect 56526 800 56634 856
rect 56802 800 56818 856
rect 56986 800 57094 856
rect 57262 800 57278 856
rect 57446 800 57554 856
rect 57722 800 57738 856
rect 57906 800 58014 856
rect 58182 800 58198 856
rect 58366 800 58474 856
rect 58642 800 58658 856
rect 58826 800 58934 856
rect 59102 800 59118 856
rect 59286 800 59394 856
rect 59562 800 59578 856
rect 59746 800 59854 856
rect 60022 800 60038 856
rect 60206 800 60314 856
rect 60482 800 60498 856
rect 60666 800 60774 856
rect 60942 800 60958 856
rect 61126 800 61234 856
rect 61402 800 61418 856
rect 61586 800 61694 856
rect 61862 800 61878 856
rect 62046 800 62154 856
rect 62322 800 62338 856
rect 62506 800 62614 856
rect 62782 800 62798 856
rect 62966 800 63074 856
rect 63242 800 63258 856
rect 63426 800 63534 856
rect 63702 800 63718 856
rect 63886 800 63994 856
rect 64162 800 64178 856
rect 64346 800 64454 856
rect 64622 800 64638 856
rect 64806 800 64914 856
rect 65082 800 65098 856
rect 65266 800 65374 856
rect 65542 800 65558 856
rect 65726 800 65834 856
rect 66002 800 66018 856
rect 66186 800 66294 856
rect 66462 800 66478 856
rect 66646 800 66754 856
rect 66922 800 66938 856
rect 67106 800 67214 856
rect 67382 800 67398 856
rect 67566 800 67674 856
rect 67842 800 67858 856
rect 68026 800 68134 856
rect 68302 800 68318 856
rect 68486 800 68594 856
rect 68762 800 68778 856
rect 68946 800 69054 856
rect 69222 800 69238 856
rect 69406 800 69514 856
rect 69682 800 69698 856
rect 69866 800 69974 856
rect 70142 800 70158 856
rect 70326 800 70342 856
rect 70510 800 70618 856
rect 70786 800 70802 856
rect 70970 800 71078 856
rect 71246 800 71262 856
rect 71430 800 71538 856
rect 71706 800 71722 856
rect 71890 800 71998 856
rect 72166 800 72182 856
rect 72350 800 72458 856
rect 72626 800 72642 856
rect 72810 800 72918 856
rect 73086 800 73102 856
rect 73270 800 73378 856
rect 73546 800 73562 856
rect 73730 800 73838 856
rect 74006 800 74022 856
rect 74190 800 74298 856
rect 74466 800 74482 856
rect 74650 800 74758 856
rect 74926 800 74942 856
rect 75110 800 75218 856
rect 75386 800 75402 856
rect 75570 800 75678 856
rect 75846 800 75862 856
rect 76030 800 76138 856
rect 76306 800 76322 856
rect 76490 800 76598 856
rect 76766 800 76782 856
rect 76950 800 77058 856
rect 77226 800 77242 856
rect 77410 800 77518 856
rect 77686 800 77702 856
rect 77870 800 77978 856
rect 78146 800 78162 856
rect 78330 800 78438 856
rect 78606 800 78622 856
rect 78790 800 78898 856
rect 79066 800 79082 856
rect 79250 800 79358 856
rect 79526 800 79542 856
rect 79710 800 79818 856
rect 79986 800 80002 856
rect 80170 800 80278 856
rect 80446 800 80462 856
rect 80630 800 80738 856
rect 80906 800 80922 856
rect 81090 800 81198 856
rect 81366 800 81382 856
rect 81550 800 81658 856
rect 81826 800 81842 856
rect 82010 800 82118 856
rect 82286 800 82302 856
rect 82470 800 82578 856
rect 82746 800 82762 856
rect 82930 800 83038 856
rect 83206 800 83222 856
rect 83390 800 83498 856
rect 83666 800 83682 856
rect 83850 800 83958 856
rect 84126 800 84142 856
rect 84310 800 84326 856
rect 84494 800 84602 856
rect 84770 800 84786 856
rect 84954 800 85062 856
rect 85230 800 85246 856
rect 85414 800 85522 856
rect 85690 800 85706 856
rect 85874 800 85982 856
rect 86150 800 86166 856
rect 86334 800 86442 856
rect 86610 800 86626 856
rect 86794 800 86902 856
rect 87070 800 87086 856
rect 87254 800 87362 856
rect 87530 800 87546 856
rect 87714 800 87822 856
rect 87990 800 88006 856
rect 88174 800 88282 856
rect 88450 800 88466 856
rect 88634 800 88742 856
rect 88910 800 88926 856
rect 89094 800 89202 856
rect 89370 800 89386 856
rect 89554 800 89662 856
rect 89830 800 89846 856
rect 90014 800 90122 856
rect 90290 800 90306 856
rect 90474 800 90582 856
rect 90750 800 90766 856
rect 90934 800 91042 856
rect 91210 800 91226 856
rect 91394 800 91502 856
rect 91670 800 91686 856
rect 91854 800 91962 856
rect 92130 800 92146 856
rect 92314 800 92422 856
rect 92590 800 92606 856
rect 92774 800 92882 856
rect 93050 800 93066 856
rect 93234 800 93342 856
rect 93510 800 93526 856
rect 93694 800 93802 856
rect 93970 800 93986 856
rect 94154 800 94262 856
rect 94430 800 94446 856
rect 94614 800 94722 856
rect 94890 800 94906 856
rect 95074 800 95182 856
rect 95350 800 95366 856
rect 95534 800 95642 856
rect 95810 800 95826 856
rect 95994 800 96102 856
rect 96270 800 96286 856
rect 96454 800 96562 856
rect 96730 800 96746 856
rect 96914 800 97022 856
rect 97190 800 97206 856
rect 97374 800 97482 856
rect 97650 800 97666 856
rect 97834 800 97942 856
rect 98110 800 98126 856
rect 98294 800 98310 856
rect 98478 800 98586 856
rect 98754 800 98770 856
rect 98938 800 99046 856
rect 99214 800 99230 856
rect 99398 800 99506 856
rect 99674 800 99690 856
rect 99858 800 99966 856
rect 100134 800 100150 856
rect 100318 800 100426 856
rect 100594 800 100610 856
rect 100778 800 100886 856
rect 101054 800 101070 856
rect 101238 800 101346 856
rect 101514 800 101530 856
rect 101698 800 101806 856
rect 101974 800 101990 856
rect 102158 800 102266 856
rect 102434 800 102450 856
rect 102618 800 102726 856
rect 102894 800 102910 856
rect 103078 800 103186 856
rect 103354 800 103370 856
rect 103538 800 103646 856
rect 103814 800 103830 856
rect 103998 800 104106 856
rect 104274 800 104290 856
rect 104458 800 104566 856
rect 104734 800 104750 856
rect 104918 800 105026 856
rect 105194 800 105210 856
rect 105378 800 105486 856
rect 105654 800 105670 856
rect 105838 800 105946 856
rect 106114 800 106130 856
rect 106298 800 106406 856
rect 106574 800 106590 856
rect 106758 800 106866 856
rect 107034 800 107050 856
rect 107218 800 107326 856
rect 107494 800 107510 856
rect 107678 800 107786 856
rect 107954 800 107970 856
rect 108138 800 108246 856
rect 108414 800 108430 856
rect 108598 800 108706 856
rect 108874 800 108890 856
rect 109058 800 109166 856
rect 109334 800 109350 856
rect 109518 800 109626 856
rect 109794 800 109810 856
rect 109978 800 110086 856
rect 110254 800 110270 856
rect 110438 800 110546 856
rect 110714 800 110730 856
rect 110898 800 111006 856
rect 111174 800 111190 856
rect 111358 800 111466 856
rect 111634 800 111650 856
rect 111818 800 111926 856
rect 112094 800 112110 856
<< metal3 >>
rect 111510 85824 112310 85944
rect 0 57264 800 57384
rect 111510 28568 112310 28688
<< obsm3 >>
rect 800 86024 111510 112097
rect 800 85744 111430 86024
rect 800 57464 111510 85744
rect 880 57184 111510 57464
rect 800 28768 111510 57184
rect 800 28488 111430 28768
rect 800 2143 111510 28488
<< metal4 >>
rect 4208 2128 4528 112112
rect 4868 2176 5188 112064
rect 5528 2176 5848 112064
rect 6188 2176 6508 112064
rect 19568 2128 19888 112112
rect 20228 2176 20548 112064
rect 20888 2176 21208 112064
rect 21548 2176 21868 112064
rect 34928 2128 35248 112112
rect 35588 2176 35908 112064
rect 36248 2176 36568 112064
rect 36908 2176 37228 112064
rect 50288 2128 50608 112112
rect 50948 2176 51268 112064
rect 51608 2176 51928 112064
rect 52268 2176 52588 112064
rect 65648 2128 65968 112112
rect 66308 2176 66628 112064
rect 66968 2176 67288 112064
rect 67628 2176 67948 112064
rect 81008 2128 81328 112112
rect 81668 2176 81988 112064
rect 82328 2176 82648 112064
rect 82988 2176 83308 112064
rect 96368 2128 96688 112112
rect 97028 2176 97348 112064
rect 97688 2176 98008 112064
rect 98348 2176 98668 112064
<< obsm4 >>
rect 16251 2619 19488 71093
rect 19968 2619 20148 71093
rect 20628 2619 20808 71093
rect 21288 2619 21468 71093
rect 21948 2619 34848 71093
rect 35328 2619 35508 71093
rect 35988 2619 36168 71093
rect 36648 2619 36828 71093
rect 37308 2619 50208 71093
rect 50688 2619 50868 71093
rect 51348 2619 51528 71093
rect 52008 2619 52188 71093
rect 52668 2619 65568 71093
rect 66048 2619 66228 71093
rect 66708 2619 66888 71093
rect 67368 2619 67548 71093
rect 68028 2619 80928 71093
rect 81408 2619 81588 71093
rect 82068 2619 82248 71093
rect 82728 2619 82908 71093
rect 83388 2619 96288 71093
rect 96768 2619 96909 71093
<< labels >>
rlabel metal2 s 478 113654 534 114454 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 30010 113654 30066 114454 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 32954 113654 33010 114454 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 35898 113654 35954 114454 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 38842 113654 38898 114454 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 41786 113654 41842 114454 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 44730 113654 44786 114454 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 47766 113654 47822 114454 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 50710 113654 50766 114454 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 53654 113654 53710 114454 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 56598 113654 56654 114454 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3422 113654 3478 114454 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 59542 113654 59598 114454 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 62486 113654 62542 114454 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 65430 113654 65486 114454 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 68466 113654 68522 114454 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 71410 113654 71466 114454 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 74354 113654 74410 114454 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 77298 113654 77354 114454 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 80242 113654 80298 114454 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 83186 113654 83242 114454 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 86130 113654 86186 114454 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6366 113654 6422 114454 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 89074 113654 89130 114454 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 92110 113654 92166 114454 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 95054 113654 95110 114454 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 97998 113654 98054 114454 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 100942 113654 100998 114454 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 103886 113654 103942 114454 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 106830 113654 106886 114454 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 109774 113654 109830 114454 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9310 113654 9366 114454 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 12254 113654 12310 114454 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 15198 113654 15254 114454 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 18142 113654 18198 114454 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 21086 113654 21142 114454 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 24122 113654 24178 114454 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 27066 113654 27122 114454 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1398 113654 1454 114454 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 31022 113654 31078 114454 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 33966 113654 34022 114454 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 36910 113654 36966 114454 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 39854 113654 39910 114454 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 42798 113654 42854 114454 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 45742 113654 45798 114454 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 48686 113654 48742 114454 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 51630 113654 51686 114454 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 54666 113654 54722 114454 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 57610 113654 57666 114454 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 4342 113654 4398 114454 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 60554 113654 60610 114454 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 63498 113654 63554 114454 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 66442 113654 66498 114454 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 69386 113654 69442 114454 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 72330 113654 72386 114454 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 75366 113654 75422 114454 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 78310 113654 78366 114454 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 81254 113654 81310 114454 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 84198 113654 84254 114454 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 87142 113654 87198 114454 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 7286 113654 7342 114454 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 90086 113654 90142 114454 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 93030 113654 93086 114454 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 95974 113654 96030 114454 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 99010 113654 99066 114454 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 101954 113654 102010 114454 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 104898 113654 104954 114454 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 107842 113654 107898 114454 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 110786 113654 110842 114454 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 10322 113654 10378 114454 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 13266 113654 13322 114454 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 16210 113654 16266 114454 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 19154 113654 19210 114454 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 22098 113654 22154 114454 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 25042 113654 25098 114454 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 27986 113654 28042 114454 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2410 113654 2466 114454 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 31942 113654 31998 114454 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 34886 113654 34942 114454 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 37922 113654 37978 114454 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 40866 113654 40922 114454 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 43810 113654 43866 114454 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 46754 113654 46810 114454 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 49698 113654 49754 114454 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 52642 113654 52698 114454 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 55586 113654 55642 114454 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 58530 113654 58586 114454 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 5354 113654 5410 114454 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 61566 113654 61622 114454 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 64510 113654 64566 114454 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 67454 113654 67510 114454 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 70398 113654 70454 114454 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 73342 113654 73398 114454 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 76286 113654 76342 114454 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 79230 113654 79286 114454 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 82174 113654 82230 114454 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 85210 113654 85266 114454 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 88154 113654 88210 114454 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 8298 113654 8354 114454 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 91098 113654 91154 114454 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 94042 113654 94098 114454 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 96986 113654 97042 114454 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 99930 113654 99986 114454 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 102874 113654 102930 114454 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 105910 113654 105966 114454 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 108854 113654 108910 114454 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 111798 113654 111854 114454 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 11242 113654 11298 114454 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 14186 113654 14242 114454 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 17222 113654 17278 114454 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 20166 113654 20222 114454 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 23110 113654 23166 114454 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 26054 113654 26110 114454 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 28998 113654 29054 114454 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 111510 28568 112310 28688 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 111510 85824 112310 85944 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 0 57264 800 57384 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 100022 0 100078 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 106922 0 106978 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 96158 0 96214 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 99562 0 99618 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 101586 0 101642 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 109222 0 109278 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 58990 0 59046 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 76838 0 76894 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 79598 0 79654 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 80334 0 80390 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 87142 0 87198 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 88522 0 88578 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 99746 0 99802 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 96368 2128 96688 112112 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 112112 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 112112 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 112112 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 81008 2128 81328 112112 6 vssd1
port 612 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 112112 6 vssd1
port 613 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 112112 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 97028 2176 97348 112064 6 vccd2
port 615 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 112064 6 vccd2
port 616 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 112064 6 vccd2
port 617 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 112064 6 vccd2
port 618 nsew power bidirectional
rlabel metal4 s 81668 2176 81988 112064 6 vssd2
port 619 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 112064 6 vssd2
port 620 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 112064 6 vssd2
port 621 nsew ground bidirectional
rlabel metal4 s 97688 2176 98008 112064 6 vdda1
port 622 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 112064 6 vdda1
port 623 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 112064 6 vdda1
port 624 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 112064 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 82328 2176 82648 112064 6 vssa1
port 626 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 112064 6 vssa1
port 627 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 112064 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 98348 2176 98668 112064 6 vdda2
port 629 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 112064 6 vdda2
port 630 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 112064 6 vdda2
port 631 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 112064 6 vdda2
port 632 nsew power bidirectional
rlabel metal4 s 82988 2176 83308 112064 6 vssa2
port 633 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 112064 6 vssa2
port 634 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 112064 6 vssa2
port 635 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 112310 114454
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 22044778
string GDS_START 1115118
<< end >>

