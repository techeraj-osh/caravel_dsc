magic
tech sky130A
magscale 1 2
timestamp 1623957084
<< obsli1 >>
rect 1104 2159 104052 105009
<< obsm1 >>
rect 106 1164 105142 105040
<< metal2 >>
rect 386 106554 442 107354
rect 1214 106554 1270 107354
rect 2134 106554 2190 107354
rect 3054 106554 3110 107354
rect 3974 106554 4030 107354
rect 4894 106554 4950 107354
rect 5814 106554 5870 107354
rect 6734 106554 6790 107354
rect 7562 106554 7618 107354
rect 8482 106554 8538 107354
rect 9402 106554 9458 107354
rect 10322 106554 10378 107354
rect 11242 106554 11298 107354
rect 12162 106554 12218 107354
rect 13082 106554 13138 107354
rect 13910 106554 13966 107354
rect 14830 106554 14886 107354
rect 15750 106554 15806 107354
rect 16670 106554 16726 107354
rect 17590 106554 17646 107354
rect 18510 106554 18566 107354
rect 19430 106554 19486 107354
rect 20258 106554 20314 107354
rect 21178 106554 21234 107354
rect 22098 106554 22154 107354
rect 23018 106554 23074 107354
rect 23938 106554 23994 107354
rect 24858 106554 24914 107354
rect 25778 106554 25834 107354
rect 26698 106554 26754 107354
rect 27526 106554 27582 107354
rect 28446 106554 28502 107354
rect 29366 106554 29422 107354
rect 30286 106554 30342 107354
rect 31206 106554 31262 107354
rect 32126 106554 32182 107354
rect 33046 106554 33102 107354
rect 33874 106554 33930 107354
rect 34794 106554 34850 107354
rect 35714 106554 35770 107354
rect 36634 106554 36690 107354
rect 37554 106554 37610 107354
rect 38474 106554 38530 107354
rect 39394 106554 39450 107354
rect 40222 106554 40278 107354
rect 41142 106554 41198 107354
rect 42062 106554 42118 107354
rect 42982 106554 43038 107354
rect 43902 106554 43958 107354
rect 44822 106554 44878 107354
rect 45742 106554 45798 107354
rect 46570 106554 46626 107354
rect 47490 106554 47546 107354
rect 48410 106554 48466 107354
rect 49330 106554 49386 107354
rect 50250 106554 50306 107354
rect 51170 106554 51226 107354
rect 52090 106554 52146 107354
rect 53010 106554 53066 107354
rect 53838 106554 53894 107354
rect 54758 106554 54814 107354
rect 55678 106554 55734 107354
rect 56598 106554 56654 107354
rect 57518 106554 57574 107354
rect 58438 106554 58494 107354
rect 59358 106554 59414 107354
rect 60186 106554 60242 107354
rect 61106 106554 61162 107354
rect 62026 106554 62082 107354
rect 62946 106554 63002 107354
rect 63866 106554 63922 107354
rect 64786 106554 64842 107354
rect 65706 106554 65762 107354
rect 66534 106554 66590 107354
rect 67454 106554 67510 107354
rect 68374 106554 68430 107354
rect 69294 106554 69350 107354
rect 70214 106554 70270 107354
rect 71134 106554 71190 107354
rect 72054 106554 72110 107354
rect 72882 106554 72938 107354
rect 73802 106554 73858 107354
rect 74722 106554 74778 107354
rect 75642 106554 75698 107354
rect 76562 106554 76618 107354
rect 77482 106554 77538 107354
rect 78402 106554 78458 107354
rect 79322 106554 79378 107354
rect 80150 106554 80206 107354
rect 81070 106554 81126 107354
rect 81990 106554 82046 107354
rect 82910 106554 82966 107354
rect 83830 106554 83886 107354
rect 84750 106554 84806 107354
rect 85670 106554 85726 107354
rect 86498 106554 86554 107354
rect 87418 106554 87474 107354
rect 88338 106554 88394 107354
rect 89258 106554 89314 107354
rect 90178 106554 90234 107354
rect 91098 106554 91154 107354
rect 92018 106554 92074 107354
rect 92846 106554 92902 107354
rect 93766 106554 93822 107354
rect 94686 106554 94742 107354
rect 95606 106554 95662 107354
rect 96526 106554 96582 107354
rect 97446 106554 97502 107354
rect 98366 106554 98422 107354
rect 99194 106554 99250 107354
rect 100114 106554 100170 107354
rect 101034 106554 101090 107354
rect 101954 106554 102010 107354
rect 102874 106554 102930 107354
rect 103794 106554 103850 107354
rect 104714 106554 104770 107354
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 754 0 810 800
rect 938 0 994 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1582 0 1638 800
rect 1766 0 1822 800
rect 2042 0 2098 800
rect 2226 0 2282 800
rect 2410 0 2466 800
rect 2686 0 2742 800
rect 2870 0 2926 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 4986 0 5042 800
rect 5262 0 5318 800
rect 5446 0 5502 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6274 0 6330 800
rect 6550 0 6606 800
rect 6734 0 6790 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8206 0 8262 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9310 0 9366 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10138 0 10194 800
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 14002 0 14058 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14646 0 14702 800
rect 14922 0 14978 800
rect 15106 0 15162 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16854 0 16910 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17682 0 17738 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18786 0 18842 800
rect 18970 0 19026 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20442 0 20498 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21730 0 21786 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24306 0 24362 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31666 0 31722 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39394 0 39450 800
rect 39578 0 39634 800
rect 39762 0 39818 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42154 0 42210 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42982 0 43038 800
rect 43258 0 43314 800
rect 43442 0 43498 800
rect 43626 0 43682 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44730 0 44786 800
rect 44914 0 44970 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48594 0 48650 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57886 0 57942 800
rect 58070 0 58126 800
rect 58254 0 58310 800
rect 58530 0 58586 800
rect 58714 0 58770 800
rect 58898 0 58954 800
rect 59174 0 59230 800
rect 59358 0 59414 800
rect 59542 0 59598 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60830 0 60886 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61474 0 61530 800
rect 61750 0 61806 800
rect 61934 0 61990 800
rect 62118 0 62174 800
rect 62394 0 62450 800
rect 62578 0 62634 800
rect 62762 0 62818 800
rect 63038 0 63094 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63682 0 63738 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64326 0 64382 800
rect 64510 0 64566 800
rect 64694 0 64750 800
rect 64970 0 65026 800
rect 65154 0 65210 800
rect 65338 0 65394 800
rect 65614 0 65670 800
rect 65798 0 65854 800
rect 65982 0 66038 800
rect 66258 0 66314 800
rect 66442 0 66498 800
rect 66626 0 66682 800
rect 66902 0 66958 800
rect 67086 0 67142 800
rect 67270 0 67326 800
rect 67546 0 67602 800
rect 67730 0 67786 800
rect 67914 0 67970 800
rect 68190 0 68246 800
rect 68374 0 68430 800
rect 68558 0 68614 800
rect 68834 0 68890 800
rect 69018 0 69074 800
rect 69202 0 69258 800
rect 69478 0 69534 800
rect 69662 0 69718 800
rect 69846 0 69902 800
rect 70122 0 70178 800
rect 70306 0 70362 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 70950 0 71006 800
rect 71134 0 71190 800
rect 71410 0 71466 800
rect 71594 0 71650 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72238 0 72294 800
rect 72422 0 72478 800
rect 72698 0 72754 800
rect 72882 0 72938 800
rect 73066 0 73122 800
rect 73342 0 73398 800
rect 73526 0 73582 800
rect 73710 0 73766 800
rect 73986 0 74042 800
rect 74170 0 74226 800
rect 74354 0 74410 800
rect 74630 0 74686 800
rect 74814 0 74870 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75458 0 75514 800
rect 75642 0 75698 800
rect 75918 0 75974 800
rect 76102 0 76158 800
rect 76286 0 76342 800
rect 76562 0 76618 800
rect 76746 0 76802 800
rect 76930 0 76986 800
rect 77206 0 77262 800
rect 77390 0 77446 800
rect 77574 0 77630 800
rect 77850 0 77906 800
rect 78034 0 78090 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78678 0 78734 800
rect 78862 0 78918 800
rect 79138 0 79194 800
rect 79322 0 79378 800
rect 79506 0 79562 800
rect 79782 0 79838 800
rect 79966 0 80022 800
rect 80150 0 80206 800
rect 80426 0 80482 800
rect 80610 0 80666 800
rect 80794 0 80850 800
rect 81070 0 81126 800
rect 81254 0 81310 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 81898 0 81954 800
rect 82082 0 82138 800
rect 82358 0 82414 800
rect 82542 0 82598 800
rect 82726 0 82782 800
rect 83002 0 83058 800
rect 83186 0 83242 800
rect 83370 0 83426 800
rect 83646 0 83702 800
rect 83830 0 83886 800
rect 84014 0 84070 800
rect 84290 0 84346 800
rect 84474 0 84530 800
rect 84658 0 84714 800
rect 84934 0 84990 800
rect 85118 0 85174 800
rect 85302 0 85358 800
rect 85578 0 85634 800
rect 85762 0 85818 800
rect 85946 0 86002 800
rect 86222 0 86278 800
rect 86406 0 86462 800
rect 86590 0 86646 800
rect 86866 0 86922 800
rect 87050 0 87106 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87694 0 87750 800
rect 87878 0 87934 800
rect 88154 0 88210 800
rect 88338 0 88394 800
rect 88522 0 88578 800
rect 88798 0 88854 800
rect 88982 0 89038 800
rect 89166 0 89222 800
rect 89442 0 89498 800
rect 89626 0 89682 800
rect 89810 0 89866 800
rect 90086 0 90142 800
rect 90270 0 90326 800
rect 90454 0 90510 800
rect 90730 0 90786 800
rect 90914 0 90970 800
rect 91098 0 91154 800
rect 91374 0 91430 800
rect 91558 0 91614 800
rect 91742 0 91798 800
rect 92018 0 92074 800
rect 92202 0 92258 800
rect 92386 0 92442 800
rect 92662 0 92718 800
rect 92846 0 92902 800
rect 93030 0 93086 800
rect 93306 0 93362 800
rect 93490 0 93546 800
rect 93674 0 93730 800
rect 93950 0 94006 800
rect 94134 0 94190 800
rect 94318 0 94374 800
rect 94594 0 94650 800
rect 94778 0 94834 800
rect 94962 0 95018 800
rect 95238 0 95294 800
rect 95422 0 95478 800
rect 95606 0 95662 800
rect 95882 0 95938 800
rect 96066 0 96122 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96710 0 96766 800
rect 96894 0 96950 800
rect 97170 0 97226 800
rect 97354 0 97410 800
rect 97538 0 97594 800
rect 97814 0 97870 800
rect 97998 0 98054 800
rect 98182 0 98238 800
rect 98458 0 98514 800
rect 98642 0 98698 800
rect 98826 0 98882 800
rect 99102 0 99158 800
rect 99286 0 99342 800
rect 99470 0 99526 800
rect 99746 0 99802 800
rect 99930 0 99986 800
rect 100114 0 100170 800
rect 100390 0 100446 800
rect 100574 0 100630 800
rect 100758 0 100814 800
rect 101034 0 101090 800
rect 101218 0 101274 800
rect 101402 0 101458 800
rect 101678 0 101734 800
rect 101862 0 101918 800
rect 102046 0 102102 800
rect 102322 0 102378 800
rect 102506 0 102562 800
rect 102690 0 102746 800
rect 102966 0 103022 800
rect 103150 0 103206 800
rect 103334 0 103390 800
rect 103610 0 103666 800
rect 103794 0 103850 800
rect 103978 0 104034 800
rect 104254 0 104310 800
rect 104438 0 104494 800
rect 104622 0 104678 800
rect 104898 0 104954 800
rect 105082 0 105138 800
<< obsm2 >>
rect 112 106498 330 106554
rect 498 106498 1158 106554
rect 1326 106498 2078 106554
rect 2246 106498 2998 106554
rect 3166 106498 3918 106554
rect 4086 106498 4838 106554
rect 5006 106498 5758 106554
rect 5926 106498 6678 106554
rect 6846 106498 7506 106554
rect 7674 106498 8426 106554
rect 8594 106498 9346 106554
rect 9514 106498 10266 106554
rect 10434 106498 11186 106554
rect 11354 106498 12106 106554
rect 12274 106498 13026 106554
rect 13194 106498 13854 106554
rect 14022 106498 14774 106554
rect 14942 106498 15694 106554
rect 15862 106498 16614 106554
rect 16782 106498 17534 106554
rect 17702 106498 18454 106554
rect 18622 106498 19374 106554
rect 19542 106498 20202 106554
rect 20370 106498 21122 106554
rect 21290 106498 22042 106554
rect 22210 106498 22962 106554
rect 23130 106498 23882 106554
rect 24050 106498 24802 106554
rect 24970 106498 25722 106554
rect 25890 106498 26642 106554
rect 26810 106498 27470 106554
rect 27638 106498 28390 106554
rect 28558 106498 29310 106554
rect 29478 106498 30230 106554
rect 30398 106498 31150 106554
rect 31318 106498 32070 106554
rect 32238 106498 32990 106554
rect 33158 106498 33818 106554
rect 33986 106498 34738 106554
rect 34906 106498 35658 106554
rect 35826 106498 36578 106554
rect 36746 106498 37498 106554
rect 37666 106498 38418 106554
rect 38586 106498 39338 106554
rect 39506 106498 40166 106554
rect 40334 106498 41086 106554
rect 41254 106498 42006 106554
rect 42174 106498 42926 106554
rect 43094 106498 43846 106554
rect 44014 106498 44766 106554
rect 44934 106498 45686 106554
rect 45854 106498 46514 106554
rect 46682 106498 47434 106554
rect 47602 106498 48354 106554
rect 48522 106498 49274 106554
rect 49442 106498 50194 106554
rect 50362 106498 51114 106554
rect 51282 106498 52034 106554
rect 52202 106498 52954 106554
rect 53122 106498 53782 106554
rect 53950 106498 54702 106554
rect 54870 106498 55622 106554
rect 55790 106498 56542 106554
rect 56710 106498 57462 106554
rect 57630 106498 58382 106554
rect 58550 106498 59302 106554
rect 59470 106498 60130 106554
rect 60298 106498 61050 106554
rect 61218 106498 61970 106554
rect 62138 106498 62890 106554
rect 63058 106498 63810 106554
rect 63978 106498 64730 106554
rect 64898 106498 65650 106554
rect 65818 106498 66478 106554
rect 66646 106498 67398 106554
rect 67566 106498 68318 106554
rect 68486 106498 69238 106554
rect 69406 106498 70158 106554
rect 70326 106498 71078 106554
rect 71246 106498 71998 106554
rect 72166 106498 72826 106554
rect 72994 106498 73746 106554
rect 73914 106498 74666 106554
rect 74834 106498 75586 106554
rect 75754 106498 76506 106554
rect 76674 106498 77426 106554
rect 77594 106498 78346 106554
rect 78514 106498 79266 106554
rect 79434 106498 80094 106554
rect 80262 106498 81014 106554
rect 81182 106498 81934 106554
rect 82102 106498 82854 106554
rect 83022 106498 83774 106554
rect 83942 106498 84694 106554
rect 84862 106498 85614 106554
rect 85782 106498 86442 106554
rect 86610 106498 87362 106554
rect 87530 106498 88282 106554
rect 88450 106498 89202 106554
rect 89370 106498 90122 106554
rect 90290 106498 91042 106554
rect 91210 106498 91962 106554
rect 92130 106498 92790 106554
rect 92958 106498 93710 106554
rect 93878 106498 94630 106554
rect 94798 106498 95550 106554
rect 95718 106498 96470 106554
rect 96638 106498 97390 106554
rect 97558 106498 98310 106554
rect 98478 106498 99138 106554
rect 99306 106498 100058 106554
rect 100226 106498 100978 106554
rect 101146 106498 101898 106554
rect 102066 106498 102818 106554
rect 102986 106498 103738 106554
rect 103906 106498 104658 106554
rect 104826 106498 105136 106554
rect 112 856 105136 106498
rect 222 800 238 856
rect 406 800 422 856
rect 590 800 698 856
rect 866 800 882 856
rect 1050 800 1066 856
rect 1234 800 1342 856
rect 1510 800 1526 856
rect 1694 800 1710 856
rect 1878 800 1986 856
rect 2154 800 2170 856
rect 2338 800 2354 856
rect 2522 800 2630 856
rect 2798 800 2814 856
rect 2982 800 2998 856
rect 3166 800 3274 856
rect 3442 800 3458 856
rect 3626 800 3642 856
rect 3810 800 3918 856
rect 4086 800 4102 856
rect 4270 800 4286 856
rect 4454 800 4562 856
rect 4730 800 4746 856
rect 4914 800 4930 856
rect 5098 800 5206 856
rect 5374 800 5390 856
rect 5558 800 5574 856
rect 5742 800 5850 856
rect 6018 800 6034 856
rect 6202 800 6218 856
rect 6386 800 6494 856
rect 6662 800 6678 856
rect 6846 800 6862 856
rect 7030 800 7138 856
rect 7306 800 7322 856
rect 7490 800 7506 856
rect 7674 800 7782 856
rect 7950 800 7966 856
rect 8134 800 8150 856
rect 8318 800 8426 856
rect 8594 800 8610 856
rect 8778 800 8794 856
rect 8962 800 9070 856
rect 9238 800 9254 856
rect 9422 800 9438 856
rect 9606 800 9714 856
rect 9882 800 9898 856
rect 10066 800 10082 856
rect 10250 800 10358 856
rect 10526 800 10542 856
rect 10710 800 10726 856
rect 10894 800 11002 856
rect 11170 800 11186 856
rect 11354 800 11370 856
rect 11538 800 11646 856
rect 11814 800 11830 856
rect 11998 800 12014 856
rect 12182 800 12290 856
rect 12458 800 12474 856
rect 12642 800 12658 856
rect 12826 800 12934 856
rect 13102 800 13118 856
rect 13286 800 13302 856
rect 13470 800 13578 856
rect 13746 800 13762 856
rect 13930 800 13946 856
rect 14114 800 14222 856
rect 14390 800 14406 856
rect 14574 800 14590 856
rect 14758 800 14866 856
rect 15034 800 15050 856
rect 15218 800 15234 856
rect 15402 800 15510 856
rect 15678 800 15694 856
rect 15862 800 15878 856
rect 16046 800 16154 856
rect 16322 800 16338 856
rect 16506 800 16522 856
rect 16690 800 16798 856
rect 16966 800 16982 856
rect 17150 800 17166 856
rect 17334 800 17442 856
rect 17610 800 17626 856
rect 17794 800 17810 856
rect 17978 800 18086 856
rect 18254 800 18270 856
rect 18438 800 18454 856
rect 18622 800 18730 856
rect 18898 800 18914 856
rect 19082 800 19098 856
rect 19266 800 19374 856
rect 19542 800 19558 856
rect 19726 800 19742 856
rect 19910 800 20018 856
rect 20186 800 20202 856
rect 20370 800 20386 856
rect 20554 800 20662 856
rect 20830 800 20846 856
rect 21014 800 21030 856
rect 21198 800 21306 856
rect 21474 800 21490 856
rect 21658 800 21674 856
rect 21842 800 21950 856
rect 22118 800 22134 856
rect 22302 800 22318 856
rect 22486 800 22594 856
rect 22762 800 22778 856
rect 22946 800 22962 856
rect 23130 800 23238 856
rect 23406 800 23422 856
rect 23590 800 23606 856
rect 23774 800 23882 856
rect 24050 800 24066 856
rect 24234 800 24250 856
rect 24418 800 24526 856
rect 24694 800 24710 856
rect 24878 800 24894 856
rect 25062 800 25170 856
rect 25338 800 25354 856
rect 25522 800 25538 856
rect 25706 800 25814 856
rect 25982 800 25998 856
rect 26166 800 26182 856
rect 26350 800 26458 856
rect 26626 800 26642 856
rect 26810 800 26826 856
rect 26994 800 27102 856
rect 27270 800 27286 856
rect 27454 800 27470 856
rect 27638 800 27746 856
rect 27914 800 27930 856
rect 28098 800 28114 856
rect 28282 800 28390 856
rect 28558 800 28574 856
rect 28742 800 28758 856
rect 28926 800 29034 856
rect 29202 800 29218 856
rect 29386 800 29402 856
rect 29570 800 29678 856
rect 29846 800 29862 856
rect 30030 800 30046 856
rect 30214 800 30322 856
rect 30490 800 30506 856
rect 30674 800 30690 856
rect 30858 800 30966 856
rect 31134 800 31150 856
rect 31318 800 31334 856
rect 31502 800 31610 856
rect 31778 800 31794 856
rect 31962 800 31978 856
rect 32146 800 32254 856
rect 32422 800 32438 856
rect 32606 800 32622 856
rect 32790 800 32898 856
rect 33066 800 33082 856
rect 33250 800 33266 856
rect 33434 800 33542 856
rect 33710 800 33726 856
rect 33894 800 33910 856
rect 34078 800 34186 856
rect 34354 800 34370 856
rect 34538 800 34554 856
rect 34722 800 34830 856
rect 34998 800 35014 856
rect 35182 800 35198 856
rect 35366 800 35474 856
rect 35642 800 35658 856
rect 35826 800 35842 856
rect 36010 800 36118 856
rect 36286 800 36302 856
rect 36470 800 36486 856
rect 36654 800 36762 856
rect 36930 800 36946 856
rect 37114 800 37130 856
rect 37298 800 37406 856
rect 37574 800 37590 856
rect 37758 800 37774 856
rect 37942 800 38050 856
rect 38218 800 38234 856
rect 38402 800 38418 856
rect 38586 800 38694 856
rect 38862 800 38878 856
rect 39046 800 39062 856
rect 39230 800 39338 856
rect 39506 800 39522 856
rect 39690 800 39706 856
rect 39874 800 39982 856
rect 40150 800 40166 856
rect 40334 800 40350 856
rect 40518 800 40626 856
rect 40794 800 40810 856
rect 40978 800 40994 856
rect 41162 800 41270 856
rect 41438 800 41454 856
rect 41622 800 41638 856
rect 41806 800 41914 856
rect 42082 800 42098 856
rect 42266 800 42282 856
rect 42450 800 42558 856
rect 42726 800 42742 856
rect 42910 800 42926 856
rect 43094 800 43202 856
rect 43370 800 43386 856
rect 43554 800 43570 856
rect 43738 800 43846 856
rect 44014 800 44030 856
rect 44198 800 44214 856
rect 44382 800 44490 856
rect 44658 800 44674 856
rect 44842 800 44858 856
rect 45026 800 45134 856
rect 45302 800 45318 856
rect 45486 800 45502 856
rect 45670 800 45778 856
rect 45946 800 45962 856
rect 46130 800 46146 856
rect 46314 800 46422 856
rect 46590 800 46606 856
rect 46774 800 46790 856
rect 46958 800 47066 856
rect 47234 800 47250 856
rect 47418 800 47434 856
rect 47602 800 47710 856
rect 47878 800 47894 856
rect 48062 800 48078 856
rect 48246 800 48354 856
rect 48522 800 48538 856
rect 48706 800 48722 856
rect 48890 800 48998 856
rect 49166 800 49182 856
rect 49350 800 49366 856
rect 49534 800 49642 856
rect 49810 800 49826 856
rect 49994 800 50010 856
rect 50178 800 50286 856
rect 50454 800 50470 856
rect 50638 800 50654 856
rect 50822 800 50930 856
rect 51098 800 51114 856
rect 51282 800 51298 856
rect 51466 800 51574 856
rect 51742 800 51758 856
rect 51926 800 51942 856
rect 52110 800 52218 856
rect 52386 800 52402 856
rect 52570 800 52678 856
rect 52846 800 52862 856
rect 53030 800 53046 856
rect 53214 800 53322 856
rect 53490 800 53506 856
rect 53674 800 53690 856
rect 53858 800 53966 856
rect 54134 800 54150 856
rect 54318 800 54334 856
rect 54502 800 54610 856
rect 54778 800 54794 856
rect 54962 800 54978 856
rect 55146 800 55254 856
rect 55422 800 55438 856
rect 55606 800 55622 856
rect 55790 800 55898 856
rect 56066 800 56082 856
rect 56250 800 56266 856
rect 56434 800 56542 856
rect 56710 800 56726 856
rect 56894 800 56910 856
rect 57078 800 57186 856
rect 57354 800 57370 856
rect 57538 800 57554 856
rect 57722 800 57830 856
rect 57998 800 58014 856
rect 58182 800 58198 856
rect 58366 800 58474 856
rect 58642 800 58658 856
rect 58826 800 58842 856
rect 59010 800 59118 856
rect 59286 800 59302 856
rect 59470 800 59486 856
rect 59654 800 59762 856
rect 59930 800 59946 856
rect 60114 800 60130 856
rect 60298 800 60406 856
rect 60574 800 60590 856
rect 60758 800 60774 856
rect 60942 800 61050 856
rect 61218 800 61234 856
rect 61402 800 61418 856
rect 61586 800 61694 856
rect 61862 800 61878 856
rect 62046 800 62062 856
rect 62230 800 62338 856
rect 62506 800 62522 856
rect 62690 800 62706 856
rect 62874 800 62982 856
rect 63150 800 63166 856
rect 63334 800 63350 856
rect 63518 800 63626 856
rect 63794 800 63810 856
rect 63978 800 63994 856
rect 64162 800 64270 856
rect 64438 800 64454 856
rect 64622 800 64638 856
rect 64806 800 64914 856
rect 65082 800 65098 856
rect 65266 800 65282 856
rect 65450 800 65558 856
rect 65726 800 65742 856
rect 65910 800 65926 856
rect 66094 800 66202 856
rect 66370 800 66386 856
rect 66554 800 66570 856
rect 66738 800 66846 856
rect 67014 800 67030 856
rect 67198 800 67214 856
rect 67382 800 67490 856
rect 67658 800 67674 856
rect 67842 800 67858 856
rect 68026 800 68134 856
rect 68302 800 68318 856
rect 68486 800 68502 856
rect 68670 800 68778 856
rect 68946 800 68962 856
rect 69130 800 69146 856
rect 69314 800 69422 856
rect 69590 800 69606 856
rect 69774 800 69790 856
rect 69958 800 70066 856
rect 70234 800 70250 856
rect 70418 800 70434 856
rect 70602 800 70710 856
rect 70878 800 70894 856
rect 71062 800 71078 856
rect 71246 800 71354 856
rect 71522 800 71538 856
rect 71706 800 71722 856
rect 71890 800 71998 856
rect 72166 800 72182 856
rect 72350 800 72366 856
rect 72534 800 72642 856
rect 72810 800 72826 856
rect 72994 800 73010 856
rect 73178 800 73286 856
rect 73454 800 73470 856
rect 73638 800 73654 856
rect 73822 800 73930 856
rect 74098 800 74114 856
rect 74282 800 74298 856
rect 74466 800 74574 856
rect 74742 800 74758 856
rect 74926 800 74942 856
rect 75110 800 75218 856
rect 75386 800 75402 856
rect 75570 800 75586 856
rect 75754 800 75862 856
rect 76030 800 76046 856
rect 76214 800 76230 856
rect 76398 800 76506 856
rect 76674 800 76690 856
rect 76858 800 76874 856
rect 77042 800 77150 856
rect 77318 800 77334 856
rect 77502 800 77518 856
rect 77686 800 77794 856
rect 77962 800 77978 856
rect 78146 800 78162 856
rect 78330 800 78438 856
rect 78606 800 78622 856
rect 78790 800 78806 856
rect 78974 800 79082 856
rect 79250 800 79266 856
rect 79434 800 79450 856
rect 79618 800 79726 856
rect 79894 800 79910 856
rect 80078 800 80094 856
rect 80262 800 80370 856
rect 80538 800 80554 856
rect 80722 800 80738 856
rect 80906 800 81014 856
rect 81182 800 81198 856
rect 81366 800 81382 856
rect 81550 800 81658 856
rect 81826 800 81842 856
rect 82010 800 82026 856
rect 82194 800 82302 856
rect 82470 800 82486 856
rect 82654 800 82670 856
rect 82838 800 82946 856
rect 83114 800 83130 856
rect 83298 800 83314 856
rect 83482 800 83590 856
rect 83758 800 83774 856
rect 83942 800 83958 856
rect 84126 800 84234 856
rect 84402 800 84418 856
rect 84586 800 84602 856
rect 84770 800 84878 856
rect 85046 800 85062 856
rect 85230 800 85246 856
rect 85414 800 85522 856
rect 85690 800 85706 856
rect 85874 800 85890 856
rect 86058 800 86166 856
rect 86334 800 86350 856
rect 86518 800 86534 856
rect 86702 800 86810 856
rect 86978 800 86994 856
rect 87162 800 87178 856
rect 87346 800 87454 856
rect 87622 800 87638 856
rect 87806 800 87822 856
rect 87990 800 88098 856
rect 88266 800 88282 856
rect 88450 800 88466 856
rect 88634 800 88742 856
rect 88910 800 88926 856
rect 89094 800 89110 856
rect 89278 800 89386 856
rect 89554 800 89570 856
rect 89738 800 89754 856
rect 89922 800 90030 856
rect 90198 800 90214 856
rect 90382 800 90398 856
rect 90566 800 90674 856
rect 90842 800 90858 856
rect 91026 800 91042 856
rect 91210 800 91318 856
rect 91486 800 91502 856
rect 91670 800 91686 856
rect 91854 800 91962 856
rect 92130 800 92146 856
rect 92314 800 92330 856
rect 92498 800 92606 856
rect 92774 800 92790 856
rect 92958 800 92974 856
rect 93142 800 93250 856
rect 93418 800 93434 856
rect 93602 800 93618 856
rect 93786 800 93894 856
rect 94062 800 94078 856
rect 94246 800 94262 856
rect 94430 800 94538 856
rect 94706 800 94722 856
rect 94890 800 94906 856
rect 95074 800 95182 856
rect 95350 800 95366 856
rect 95534 800 95550 856
rect 95718 800 95826 856
rect 95994 800 96010 856
rect 96178 800 96194 856
rect 96362 800 96470 856
rect 96638 800 96654 856
rect 96822 800 96838 856
rect 97006 800 97114 856
rect 97282 800 97298 856
rect 97466 800 97482 856
rect 97650 800 97758 856
rect 97926 800 97942 856
rect 98110 800 98126 856
rect 98294 800 98402 856
rect 98570 800 98586 856
rect 98754 800 98770 856
rect 98938 800 99046 856
rect 99214 800 99230 856
rect 99398 800 99414 856
rect 99582 800 99690 856
rect 99858 800 99874 856
rect 100042 800 100058 856
rect 100226 800 100334 856
rect 100502 800 100518 856
rect 100686 800 100702 856
rect 100870 800 100978 856
rect 101146 800 101162 856
rect 101330 800 101346 856
rect 101514 800 101622 856
rect 101790 800 101806 856
rect 101974 800 101990 856
rect 102158 800 102266 856
rect 102434 800 102450 856
rect 102618 800 102634 856
rect 102802 800 102910 856
rect 103078 800 103094 856
rect 103262 800 103278 856
rect 103446 800 103554 856
rect 103722 800 103738 856
rect 103906 800 103922 856
rect 104090 800 104198 856
rect 104366 800 104382 856
rect 104550 800 104566 856
rect 104734 800 104842 856
rect 105010 800 105026 856
<< metal3 >>
rect 104410 53592 105210 53712
<< obsm3 >>
rect 2497 53792 104410 105025
rect 2497 53512 104330 53792
rect 2497 2143 104410 53512
<< metal4 >>
rect 4208 2128 4528 105040
rect 4868 2176 5188 104992
rect 5528 2176 5848 104992
rect 6188 2176 6508 104992
rect 19568 2128 19888 105040
rect 20228 2176 20548 104992
rect 20888 2176 21208 104992
rect 21548 2176 21868 104992
rect 34928 2128 35248 105040
rect 35588 2176 35908 104992
rect 36248 2176 36568 104992
rect 36908 2176 37228 104992
rect 50288 2128 50608 105040
rect 50948 2176 51268 104992
rect 51608 2176 51928 104992
rect 52268 2176 52588 104992
rect 65648 2128 65968 105040
rect 66308 2176 66628 104992
rect 66968 2176 67288 104992
rect 67628 2176 67948 104992
rect 81008 2128 81328 105040
rect 81668 2176 81988 104992
rect 82328 2176 82648 104992
rect 82988 2176 83308 104992
rect 96368 2128 96688 105040
rect 97028 2176 97348 104992
rect 97688 2176 98008 104992
rect 98348 2176 98668 104992
<< obsm4 >>
rect 12939 2211 19488 103597
rect 19968 2211 20148 103597
rect 20628 2211 20808 103597
rect 21288 2211 21468 103597
rect 21948 2211 34717 103597
<< labels >>
rlabel metal2 s 386 106554 442 107354 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 27526 106554 27582 107354 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 30286 106554 30342 107354 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 33046 106554 33102 107354 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 35714 106554 35770 107354 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 38474 106554 38530 107354 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 41142 106554 41198 107354 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 43902 106554 43958 107354 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 46570 106554 46626 107354 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 49330 106554 49386 107354 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 52090 106554 52146 107354 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3054 106554 3110 107354 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 54758 106554 54814 107354 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 57518 106554 57574 107354 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 60186 106554 60242 107354 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 62946 106554 63002 107354 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 65706 106554 65762 107354 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 68374 106554 68430 107354 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 71134 106554 71190 107354 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 73802 106554 73858 107354 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 76562 106554 76618 107354 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 79322 106554 79378 107354 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5814 106554 5870 107354 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 81990 106554 82046 107354 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 84750 106554 84806 107354 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 87418 106554 87474 107354 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 90178 106554 90234 107354 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 92846 106554 92902 107354 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 95606 106554 95662 107354 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 98366 106554 98422 107354 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 101034 106554 101090 107354 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 8482 106554 8538 107354 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 11242 106554 11298 107354 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 13910 106554 13966 107354 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 16670 106554 16726 107354 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 19430 106554 19486 107354 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 22098 106554 22154 107354 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 24858 106554 24914 107354 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1214 106554 1270 107354 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 28446 106554 28502 107354 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 31206 106554 31262 107354 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 33874 106554 33930 107354 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 36634 106554 36690 107354 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 39394 106554 39450 107354 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 42062 106554 42118 107354 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 44822 106554 44878 107354 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 47490 106554 47546 107354 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 50250 106554 50306 107354 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 53010 106554 53066 107354 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3974 106554 4030 107354 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 55678 106554 55734 107354 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 58438 106554 58494 107354 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 61106 106554 61162 107354 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 63866 106554 63922 107354 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 66534 106554 66590 107354 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 69294 106554 69350 107354 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 72054 106554 72110 107354 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 74722 106554 74778 107354 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 77482 106554 77538 107354 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 80150 106554 80206 107354 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6734 106554 6790 107354 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 82910 106554 82966 107354 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 85670 106554 85726 107354 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 88338 106554 88394 107354 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 91098 106554 91154 107354 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 93766 106554 93822 107354 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 96526 106554 96582 107354 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 99194 106554 99250 107354 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 101954 106554 102010 107354 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 9402 106554 9458 107354 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 12162 106554 12218 107354 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 14830 106554 14886 107354 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 17590 106554 17646 107354 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 20258 106554 20314 107354 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 23018 106554 23074 107354 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 25778 106554 25834 107354 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2134 106554 2190 107354 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 29366 106554 29422 107354 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 32126 106554 32182 107354 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 34794 106554 34850 107354 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 37554 106554 37610 107354 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 40222 106554 40278 107354 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 42982 106554 43038 107354 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 45742 106554 45798 107354 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 48410 106554 48466 107354 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 51170 106554 51226 107354 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 53838 106554 53894 107354 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4894 106554 4950 107354 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 56598 106554 56654 107354 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 59358 106554 59414 107354 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 62026 106554 62082 107354 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 64786 106554 64842 107354 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 67454 106554 67510 107354 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 70214 106554 70270 107354 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 72882 106554 72938 107354 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 75642 106554 75698 107354 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 78402 106554 78458 107354 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 81070 106554 81126 107354 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 7562 106554 7618 107354 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 83830 106554 83886 107354 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 86498 106554 86554 107354 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 89258 106554 89314 107354 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 92018 106554 92074 107354 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 94686 106554 94742 107354 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 97446 106554 97502 107354 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 100114 106554 100170 107354 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 102874 106554 102930 107354 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 10322 106554 10378 107354 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 13082 106554 13138 107354 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 15750 106554 15806 107354 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 18510 106554 18566 107354 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 21178 106554 21234 107354 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 23938 106554 23994 107354 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 26698 106554 26754 107354 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 103794 106554 103850 107354 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 104410 53592 105210 53712 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 104714 106554 104770 107354 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 79506 0 79562 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 87510 0 87566 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 94594 0 94650 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 99746 0 99802 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 61106 0 61162 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 64970 0 65026 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 66902 0 66958 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 67546 0 67602 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 81714 0 81770 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 84290 0 84346 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 294 0 350 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 754 0 810 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 22650 0 22706 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 96368 2128 96688 105040 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 105040 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 105040 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 105040 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 81008 2128 81328 105040 6 vssd1
port 612 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 105040 6 vssd1
port 613 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 105040 6 vssd1
port 614 nsew ground bidirectional
rlabel metal4 s 97028 2176 97348 104992 6 vccd2
port 615 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 104992 6 vccd2
port 616 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 104992 6 vccd2
port 617 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 104992 6 vccd2
port 618 nsew power bidirectional
rlabel metal4 s 81668 2176 81988 104992 6 vssd2
port 619 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 104992 6 vssd2
port 620 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 104992 6 vssd2
port 621 nsew ground bidirectional
rlabel metal4 s 97688 2176 98008 104992 6 vdda1
port 622 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 104992 6 vdda1
port 623 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 104992 6 vdda1
port 624 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 104992 6 vdda1
port 625 nsew power bidirectional
rlabel metal4 s 82328 2176 82648 104992 6 vssa1
port 626 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 104992 6 vssa1
port 627 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 104992 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 98348 2176 98668 104992 6 vdda2
port 629 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 104992 6 vdda2
port 630 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 104992 6 vdda2
port 631 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 104992 6 vdda2
port 632 nsew power bidirectional
rlabel metal4 s 82988 2176 83308 104992 6 vssa2
port 633 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 104992 6 vssa2
port 634 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 104992 6 vssa2
port 635 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 105210 107354
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 19855326
string GDS_START 1096902
<< end >>

