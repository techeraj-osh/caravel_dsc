* NGSPICE file created from user_proj_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102]
+ la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107]
+ la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112]
+ la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122]
+ la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66]
+ la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77]
+ la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88]
+ la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3]
+ wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i
+ wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2 vdda2_uq0 vdda2_uq1
+ vdda2_uq2 vdda1_uq0 vdda1_uq1 vdda1_uq2 vccd2_uq0 vccd2_uq1 vccd2_uq2 vssa2_uq0
+ vssa2_uq1 vssa1_uq0 vssa1_uq1 vssd2_uq0 vssd2_uq1
X_09671_ _09671_/A _09671_/B vssd1 vssd1 vccd1 vccd1 _09671_/Y sky130_fd_sc_hd__nor2_1
X_06883_ _06883_/A _06883_/B vssd1 vssd1 vccd1 vccd1 _06883_/Y sky130_fd_sc_hd__nor2_1
X_08622_ _11941_/X _08608_/X _12732_/Q _08610_/X vssd1 vssd1 vccd1 vccd1 _12732_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08553_ _12751_/Q vssd1 vssd1 vccd1 vccd1 _08553_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07504_ _13007_/Q vssd1 vssd1 vccd1 vccd1 _09284_/C sky130_fd_sc_hd__inv_2
X_08484_ _08471_/Y _07821_/X _13042_/Q _07822_/Y _08483_/X vssd1 vssd1 vccd1 vccd1
+ _08484_/X sky130_fd_sc_hd__a221o_1
XPHY_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07435_ _07443_/A vssd1 vssd1 vccd1 vccd1 _07435_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07366_ _11432_/X _07353_/X _13056_/Q _07354_/X vssd1 vssd1 vccd1 vccd1 _13056_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09105_ _12531_/Q _09099_/X input342/X _09100_/X vssd1 vssd1 vccd1 vccd1 _12531_/D
+ sky130_fd_sc_hd__a22o_1
X_06317_ _06303_/X _06314_/X _06316_/X _13262_/Q _06306_/X vssd1 vssd1 vccd1 vccd1
+ _13262_/D sky130_fd_sc_hd__a32o_1
X_07297_ _13078_/Q _07285_/X _07296_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _13078_/D
+ sky130_fd_sc_hd__a22o_1
X_09036_ _09283_/A _09036_/B vssd1 vssd1 vccd1 vccd1 _12572_/D sky130_fd_sc_hd__nor2_1
X_06248_ _06241_/Y _06196_/X _06241_/Y _06196_/X vssd1 vssd1 vccd1 vccd1 _06248_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_163_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06179_ _06179_/A vssd1 vssd1 vccd1 vccd1 _06179_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09938_ _09949_/A vssd1 vssd1 vccd1 vccd1 _09938_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09869_ _09880_/A _09867_/X _09785_/A _09868_/X _09857_/Y vssd1 vssd1 vccd1 vccd1
+ _09871_/B sky130_fd_sc_hd__o221a_1
XFILLER_46_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11900_ _10740_/X _10743_/X _12193_/S vssd1 vssd1 vccd1 vccd1 _11900_/X sky130_fd_sc_hd__mux2_1
XPHY_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _12880_/CLK _12880_/D _08012_/X vssd1 vssd1 vccd1 vccd1 _12880_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _09927_/Y _12856_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11831_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11762_ _11761_/X _12104_/X _11774_/S vssd1 vssd1 vccd1 vccd1 _12430_/D sky130_fd_sc_hd__mux2_1
XPHY_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10713_ _13239_/Q _11111_/A _10686_/A _10788_/A _06448_/Y vssd1 vssd1 vccd1 vccd1
+ _11051_/A sky130_fd_sc_hd__o221a_1
XPHY_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11405_/X _09179_/B _11703_/S vssd1 vssd1 vccd1 vccd1 _11693_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10644_ _08929_/A _08929_/B _10643_/Y vssd1 vssd1 vccd1 vccd1 _10644_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10575_ _12399_/D _12400_/D vssd1 vssd1 vccd1 vccd1 _10579_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12314_ _12987_/CLK _12314_/D vssd1 vssd1 vccd1 vccd1 _12314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12245_ _12777_/Q _12850_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12245_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12176_ _11143_/X _11138_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _12176_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11127_ _11033_/A _10788_/X _13243_/Q _11111_/X _11112_/X vssd1 vssd1 vccd1 vccd1
+ _11127_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11058_ _11058_/A vssd1 vssd1 vccd1 vccd1 _11058_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_wb_clk_i _12960_/CLK vssd1 vssd1 vccd1 vccd1 _12586_/CLK sky130_fd_sc_hd__clkbuf_16
X_10009_ _08753_/Y _10003_/X _06195_/Y _09972_/A _09991_/A vssd1 vssd1 vccd1 vccd1
+ _10009_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07220_ _11572_/X _07218_/X _13107_/Q _07219_/X vssd1 vssd1 vccd1 vccd1 _13107_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07151_ _11532_/X _07145_/X _13131_/Q _07146_/X vssd1 vssd1 vccd1 vccd1 _13131_/D
+ sky130_fd_sc_hd__a22o_1
X_06102_ _06102_/A vssd1 vssd1 vccd1 vccd1 _06103_/B sky130_fd_sc_hd__inv_2
X_07082_ _07069_/X _07074_/X _06351_/X _13147_/Q _07042_/A vssd1 vssd1 vccd1 vccd1
+ _13147_/D sky130_fd_sc_hd__a32o_1
XFILLER_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput401 _10112_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput412 _11194_/LO vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__clkbuf_2
X_06033_ _12715_/Q vssd1 vssd1 vccd1 vccd1 _06033_/Y sky130_fd_sc_hd__inv_2
Xoutput423 _11204_/LO vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__clkbuf_2
Xoutput434 _11214_/LO vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput445 _09334_/X vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__clkbuf_2
Xoutput456 _11325_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput467 _11335_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__clkbuf_2
Xoutput478 _11229_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput489 _11239_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07984_ _12890_/Q _07974_/X _07983_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _12890_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09723_ _13208_/Q _13207_/Q _06705_/Y _06710_/Y vssd1 vssd1 vccd1 vccd1 _09725_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06935_ _06935_/A _06935_/B vssd1 vssd1 vccd1 vccd1 _06935_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09654_ _13197_/Q _09653_/A _09652_/Y _09653_/Y vssd1 vssd1 vccd1 vccd1 _09655_/B
+ sky130_fd_sc_hd__a22o_2
X_06866_ _06526_/X _06857_/B _06864_/Y _06556_/X _06865_/Y vssd1 vssd1 vccd1 vccd1
+ _06867_/A sky130_fd_sc_hd__o32a_1
X_08605_ _11947_/X _08592_/X _12738_/Q _08593_/X vssd1 vssd1 vccd1 vccd1 _12738_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06797_ _06783_/A _06783_/B _06783_/X vssd1 vssd1 vccd1 vccd1 _06797_/X sky130_fd_sc_hd__a21bo_1
X_09585_ _13156_/Q _07737_/A _09584_/Y _09478_/X vssd1 vssd1 vccd1 vccd1 _09585_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_83_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08536_ _08504_/A _12236_/X _06396_/A _10691_/B vssd1 vssd1 vccd1 vccd1 _12755_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_169_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08467_ _08467_/A _08467_/B _08467_/C _08466_/X vssd1 vssd1 vccd1 vccd1 _08474_/C
+ sky130_fd_sc_hd__or4b_4
XPHY_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07418_ _07428_/A vssd1 vssd1 vccd1 vccd1 _07418_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08398_ _09978_/B vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__buf_2
XFILLER_177_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07349_ _11439_/X _07338_/X _13063_/Q _07339_/X vssd1 vssd1 vccd1 vccd1 _13063_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10360_ _10371_/A _10360_/B _10360_/C vssd1 vssd1 vccd1 vccd1 _10360_/Y sky130_fd_sc_hd__nor3_1
XFILLER_164_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09019_ _09019_/A _09019_/B _11635_/X vssd1 vssd1 vccd1 vccd1 _12579_/D sky130_fd_sc_hd__and3_1
XFILLER_88_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10291_ _09931_/Y _09968_/X _10282_/X _10290_/X vssd1 vssd1 vccd1 vccd1 _10291_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12030_ _11088_/X _11078_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12030_/X sky130_fd_sc_hd__mux2_4
XFILLER_105_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12932_ _12973_/CLK _12932_/D vssd1 vssd1 vccd1 vccd1 _12932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _12864_/CLK _12863_/D _08057_/X vssd1 vssd1 vccd1 vccd1 _12863_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _12086_/X _11813_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11814_/X sky130_fd_sc_hd__mux2_1
XPHY_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12864_/CLK _12794_/D _08381_/X vssd1 vssd1 vccd1 vccd1 _12794_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11372_/X _11744_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11745_/X sky130_fd_sc_hd__mux2_1
XPHY_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _11675_/X _11385_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12380_/D sky130_fd_sc_hd__mux2_1
XPHY_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10627_ _10627_/A _11817_/S _10627_/C vssd1 vssd1 vccd1 vccd1 _10627_/X sky130_fd_sc_hd__and3_1
XFILLER_127_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10558_ _10558_/A _10558_/B vssd1 vssd1 vccd1 vccd1 _10558_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13277_ _13279_/CLK _13277_/D _06230_/X vssd1 vssd1 vccd1 vccd1 _13277_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10489_ _12494_/Q vssd1 vssd1 vccd1 vccd1 _10489_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12228_ _12227_/X _12634_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12228_/X sky130_fd_sc_hd__mux2_2
XFILLER_194_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12159_ _10013_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12159_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06720_ _06720_/A _06720_/B vssd1 vssd1 vccd1 vccd1 _06720_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06651_ _13214_/Q vssd1 vssd1 vccd1 vccd1 _06651_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09370_ _09363_/Y _12414_/Q _09366_/Y _12399_/Q _09369_/X vssd1 vssd1 vccd1 vccd1
+ _09371_/D sky130_fd_sc_hd__a221oi_2
X_06582_ _12759_/Q _12758_/Q vssd1 vssd1 vccd1 vccd1 _06583_/A sky130_fd_sc_hd__and2_1
XFILLER_75_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08321_ _12818_/Q _11593_/X _08321_/S vssd1 vssd1 vccd1 vccd1 _12818_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08252_ _12843_/Q _08251_/X _07287_/X _11417_/S vssd1 vssd1 vccd1 vccd1 _12843_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07203_ _07264_/A vssd1 vssd1 vccd1 vccd1 _07249_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_192_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08183_ _13136_/Q vssd1 vssd1 vccd1 vccd1 _08183_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07134_ _11539_/X _07130_/X _13138_/Q _07131_/X vssd1 vssd1 vccd1 vccd1 _13138_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07065_ _07154_/A vssd1 vssd1 vccd1 vccd1 _07078_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_160_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06016_ _12607_/Q vssd1 vssd1 vccd1 vccd1 _08556_/D sky130_fd_sc_hd__inv_2
XFILLER_160_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07967_ _12893_/Q _11482_/X _07967_/S vssd1 vssd1 vccd1 vccd1 _12893_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09706_ _09706_/A vssd1 vssd1 vccd1 vccd1 _09706_/Y sky130_fd_sc_hd__inv_2
X_06918_ _11100_/A _06918_/B vssd1 vssd1 vccd1 vccd1 _06918_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07898_ _12922_/Q _11511_/X _07904_/S vssd1 vssd1 vccd1 vccd1 _12922_/D sky130_fd_sc_hd__mux2_1
XFILLER_83_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09637_ _13194_/Q vssd1 vssd1 vccd1 vccd1 _09637_/Y sky130_fd_sc_hd__inv_2
X_06849_ _12025_/X _12021_/X _12025_/X _12021_/X vssd1 vssd1 vccd1 vccd1 _06849_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_128_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09568_ _09568_/A _09568_/B vssd1 vssd1 vccd1 vccd1 _09568_/Y sky130_fd_sc_hd__nand2_1
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ _08519_/A vssd1 vssd1 vccd1 vccd1 _08519_/X sky130_fd_sc_hd__clkbuf_2
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09499_ _13169_/Q vssd1 vssd1 vccd1 vccd1 _09500_/B sky130_fd_sc_hd__inv_2
XFILLER_130_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11530_ _12819_/Q _10528_/B _11533_/S vssd1 vssd1 vccd1 vccd1 _11530_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11461_ _12904_/Q _09244_/B _11469_/S vssd1 vssd1 vccd1 vccd1 _11461_/X sky130_fd_sc_hd__mux2_1
XPHY_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13200_ _13201_/CLK _13200_/D _06777_/X vssd1 vssd1 vccd1 vccd1 _13200_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10412_ _10412_/A _10413_/B _10474_/A vssd1 vssd1 vccd1 vccd1 _10412_/Y sky130_fd_sc_hd__nor3_2
X_11392_ _10574_/Y _12399_/D _11392_/S vssd1 vssd1 vccd1 vccd1 _11392_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13131_ _12168_/X _13131_/D _07150_/X vssd1 vssd1 vccd1 vccd1 _13131_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10343_ _10346_/C vssd1 vssd1 vccd1 vccd1 _10344_/B sky130_fd_sc_hd__inv_2
XFILLER_180_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13062_ _12165_/X _13062_/D _07350_/X vssd1 vssd1 vccd1 vccd1 _13062_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10274_ _09928_/Y _09968_/X _10265_/X _10273_/X vssd1 vssd1 vccd1 vccd1 _10274_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_79_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12013_ _11065_/X _11057_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _12013_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12915_ _12166_/X _12915_/D _07913_/X vssd1 vssd1 vccd1 vccd1 _12915_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12846_ _12868_/CLK _12846_/D _08101_/X vssd1 vssd1 vccd1 vccd1 _12846_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12779_/CLK _12777_/D _08427_/X vssd1 vssd1 vccd1 vccd1 _12777_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11728_ _09179_/A _11727_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11728_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11659_ _10522_/Y _10558_/Y _11675_/S vssd1 vssd1 vccd1 vccd1 _11659_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08870_ _07747_/X _06342_/Y _08837_/A _12640_/Q vssd1 vssd1 vccd1 vccd1 _12640_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_123_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07821_ _12901_/Q vssd1 vssd1 vccd1 vccd1 _07821_/X sky130_fd_sc_hd__buf_2
XFILLER_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07752_ _12307_/Q vssd1 vssd1 vccd1 vccd1 _07752_/Y sky130_fd_sc_hd__inv_2
X_06703_ _06700_/X _06701_/X _11989_/X _06702_/X vssd1 vssd1 vccd1 vccd1 _06703_/X
+ sky130_fd_sc_hd__o22a_1
X_07683_ _07668_/C _07648_/A _12573_/Q vssd1 vssd1 vccd1 vccd1 _07686_/A sky130_fd_sc_hd__o21a_1
XFILLER_38_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09422_ _09422_/A _09422_/B _09422_/C _09421_/X vssd1 vssd1 vccd1 vccd1 _09431_/B
+ sky130_fd_sc_hd__or4b_4
X_06634_ _06634_/A _12758_/Q vssd1 vssd1 vccd1 vccd1 _06636_/A sky130_fd_sc_hd__or2b_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09353_ _09340_/X _09353_/B _09353_/C _09353_/D vssd1 vssd1 vccd1 vccd1 _09353_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_178_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06565_ _12178_/X _12177_/X _12178_/X _12177_/X vssd1 vssd1 vccd1 vccd1 _06565_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08304_ _08311_/A vssd1 vssd1 vccd1 vccd1 _08304_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09284_ _09284_/A _09284_/B _09284_/C vssd1 vssd1 vccd1 vccd1 _09284_/X sky130_fd_sc_hd__or3_1
X_06496_ _12040_/X _06494_/Y _12040_/X _06494_/Y vssd1 vssd1 vccd1 vccd1 _06497_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_127_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08235_ _13100_/Q _10454_/B _13093_/Q _10433_/A vssd1 vssd1 vccd1 vccd1 _08237_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_197_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08166_ _13138_/Q _08164_/Y _08165_/Y _12809_/Q vssd1 vssd1 vccd1 vccd1 _08166_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07117_ _11546_/X _07113_/X _13145_/Q _07116_/X vssd1 vssd1 vccd1 vccd1 _13145_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ _12848_/Q _08082_/A _07300_/X _08083_/A vssd1 vssd1 vccd1 vccd1 _12848_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07048_ _07477_/A vssd1 vssd1 vccd1 vccd1 _07154_/A sky130_fd_sc_hd__buf_6
XFILLER_134_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08999_ _12936_/Q _12934_/Q vssd1 vssd1 vccd1 vccd1 _08999_/X sky130_fd_sc_hd__or2_1
XFILLER_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_117_wb_clk_i _12726_/CLK vssd1 vssd1 vccd1 vccd1 _12719_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10961_ _10977_/B _10960_/X _10977_/B _10960_/X vssd1 vssd1 vccd1 vccd1 _12347_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12700_ _12717_/CLK _12700_/D _08704_/X vssd1 vssd1 vccd1 vccd1 _12700_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10892_ _12524_/Q _12336_/Q _12525_/Q _12337_/Q _10891_/X vssd1 vssd1 vccd1 vccd1
+ _10892_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12631_ _13156_/CLK _12631_/D _08892_/X vssd1 vssd1 vccd1 vccd1 _12631_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12562_ _13283_/CLK _12562_/D vssd1 vssd1 vccd1 vccd1 _12562_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11513_ _10400_/X _10793_/A _11513_/S vssd1 vssd1 vccd1 vccd1 _11513_/X sky130_fd_sc_hd__mux2_1
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _12939_/CLK _12493_/D vssd1 vssd1 vccd1 vccd1 _12493_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11444_ _12919_/Q _10794_/D _11449_/S vssd1 vssd1 vccd1 vccd1 _11444_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11375_ _10665_/Y _12428_/Q _12103_/S vssd1 vssd1 vccd1 vccd1 _11375_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13114_ _12168_/X _13114_/D _07192_/X vssd1 vssd1 vccd1 vccd1 _13114_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10326_ _12896_/Q _10326_/B vssd1 vssd1 vccd1 vccd1 _10328_/B sky130_fd_sc_hd__nand2_2
XFILLER_180_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13045_ _12165_/X _13045_/D _07394_/X vssd1 vssd1 vccd1 vccd1 _13045_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10257_ _10252_/Y _10163_/X _10253_/Y _10165_/X _10256_/X vssd1 vssd1 vccd1 vccd1
+ _10257_/X sky130_fd_sc_hd__o221a_1
XFILLER_78_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10188_ _10181_/Y _10140_/X _09544_/Y _10141_/X _10187_/X vssd1 vssd1 vccd1 vccd1
+ _10188_/X sky130_fd_sc_hd__o221a_1
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12829_ _12169_/X _12829_/D _08293_/X vssd1 vssd1 vccd1 vccd1 _12829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06350_ _12944_/Q _06120_/X _12944_/Q _06120_/X vssd1 vssd1 vccd1 vccd1 _06351_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06281_ _06281_/A vssd1 vssd1 vccd1 vccd1 _06281_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08020_ _08038_/A vssd1 vssd1 vccd1 vccd1 _08036_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09971_ _09999_/A vssd1 vssd1 vccd1 vccd1 _09972_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08922_ _12419_/Q vssd1 vssd1 vccd1 vccd1 _08926_/A sky130_fd_sc_hd__inv_2
XFILLER_112_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08853_ _08849_/X _06305_/X _08852_/X _12647_/Q vssd1 vssd1 vccd1 vccd1 _12647_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07804_ _12900_/Q vssd1 vssd1 vccd1 vccd1 _07804_/X sky130_fd_sc_hd__buf_2
X_08784_ _12673_/Q vssd1 vssd1 vccd1 vccd1 _08784_/Y sky130_fd_sc_hd__inv_2
X_07735_ _07735_/A vssd1 vssd1 vccd1 vccd1 _09475_/A sky130_fd_sc_hd__inv_2
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07666_ _07666_/A vssd1 vssd1 vccd1 vccd1 _07666_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _12412_/D vssd1 vssd1 vccd1 vccd1 _10611_/B sky130_fd_sc_hd__inv_2
XFILLER_198_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06617_ _06610_/X _06614_/X _06620_/A vssd1 vssd1 vccd1 vccd1 _06625_/A sky130_fd_sc_hd__a21oi_1
X_07597_ _12574_/Q vssd1 vssd1 vccd1 vccd1 _07598_/C sky130_fd_sc_hd__inv_2
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09336_ _12452_/Q vssd1 vssd1 vccd1 vccd1 _09336_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06548_ _06548_/A vssd1 vssd1 vccd1 vccd1 _06548_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09267_ _09433_/B _09267_/B _09267_/C _09433_/A vssd1 vssd1 vccd1 vccd1 _09267_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_193_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06479_ _11885_/X _06479_/B vssd1 vssd1 vccd1 vccd1 _06479_/Y sky130_fd_sc_hd__nand2_1
XFILLER_194_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08218_ _08205_/Y _08128_/X _13109_/Q _10477_/A vssd1 vssd1 vccd1 vccd1 _08218_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_181_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09198_ _12487_/Q _09190_/X _09180_/D _09192_/X vssd1 vssd1 vccd1 vccd1 _12487_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08149_ _12818_/Q vssd1 vssd1 vccd1 vccd1 _10444_/B sky130_fd_sc_hd__inv_2
XFILLER_134_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11160_ vssd1 vssd1 vccd1 vccd1 _11160_/HI _11160_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10111_ _08197_/Y _10070_/X _10110_/X vssd1 vssd1 vccd1 vccd1 _10111_/Y sky130_fd_sc_hd__o21ai_1
X_11091_ _10767_/X _11054_/X _06383_/X _11055_/X _11060_/X vssd1 vssd1 vccd1 vccd1
+ _11091_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput301 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 _07095_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput312 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _07096_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_1_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10042_ _10190_/A vssd1 vssd1 vccd1 vccd1 _10150_/A sky130_fd_sc_hd__clkbuf_2
Xinput323 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _11967_/S sky130_fd_sc_hd__buf_4
Xinput334 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 _07980_/A sky130_fd_sc_hd__buf_2
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput345 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 _10792_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_102_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput356 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 input356/X sky130_fd_sc_hd__buf_4
XFILLER_102_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11993_ _11102_/X _11094_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _11993_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944_ _10944_/A vssd1 vssd1 vccd1 vccd1 _10944_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10875_ _10861_/Y _10862_/Y _10890_/A _10869_/X vssd1 vssd1 vccd1 vccd1 _10876_/A
+ sky130_fd_sc_hd__o22a_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _12664_/CLK _12614_/D _08964_/X vssd1 vssd1 vccd1 vccd1 _12614_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _13241_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12545_ _13001_/CLK _12545_/D vssd1 vssd1 vccd1 vccd1 _12545_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_14_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12467_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12476_ _12477_/CLK _12476_/D vssd1 vssd1 vccd1 vccd1 _12476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11427_ _12902_/Q input360/X _11433_/S vssd1 vssd1 vccd1 vccd1 _11427_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11358_ _09330_/A _10545_/Y _12321_/Q vssd1 vssd1 vccd1 vccd1 _11358_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10309_ _13023_/Q _10276_/X _13056_/Q _10277_/X vssd1 vssd1 vccd1 vccd1 _10309_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11289_ vssd1 vssd1 vccd1 vccd1 _11289_/HI _11289_/LO sky130_fd_sc_hd__conb_1
X_13028_ _12164_/X _13028_/D _07443_/X vssd1 vssd1 vccd1 vccd1 _13028_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07520_ _07520_/A vssd1 vssd1 vccd1 vccd1 _07520_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07451_ _11467_/X _07444_/X _13026_/Q _07445_/X vssd1 vssd1 vccd1 vccd1 _13026_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06402_ _06412_/A vssd1 vssd1 vccd1 vccd1 _06402_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07382_ _11426_/X _07368_/X _13050_/Q _07369_/X vssd1 vssd1 vccd1 vccd1 _13050_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09121_ _12519_/Q _09115_/X _07997_/X _09116_/X vssd1 vssd1 vccd1 vccd1 _12519_/D
+ sky130_fd_sc_hd__a22o_1
X_06333_ _06303_/X _06314_/X _06332_/Y _13259_/Q _06306_/X vssd1 vssd1 vccd1 vccd1
+ _13259_/D sky130_fd_sc_hd__a32o_1
XFILLER_176_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06264_ _06134_/Y _06069_/A _06064_/A vssd1 vssd1 vccd1 vccd1 _06264_/Y sky130_fd_sc_hd__o21ai_1
X_09052_ _10244_/A vssd1 vssd1 vccd1 vccd1 _09058_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_191_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08003_ _12884_/Q _07996_/X _07290_/X _07998_/X vssd1 vssd1 vccd1 vccd1 _12884_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06195_ _13283_/Q vssd1 vssd1 vccd1 vccd1 _06195_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ _08770_/Y _09952_/X _06228_/X _09949_/X _09950_/X vssd1 vssd1 vccd1 vccd1
+ _09954_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_44_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08905_ _08912_/A vssd1 vssd1 vccd1 vccd1 _08905_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09885_ _09686_/X _09884_/A _13238_/Q _09884_/Y _09492_/A vssd1 vssd1 vccd1 vccd1
+ _09886_/B sky130_fd_sc_hd__o221a_1
XFILLER_135_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08836_ _08836_/A vssd1 vssd1 vccd1 vccd1 _08836_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ _12678_/Q vssd1 vssd1 vccd1 vccd1 _08767_/Y sky130_fd_sc_hd__inv_2
XPHY_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07718_ _12310_/Q vssd1 vssd1 vccd1 vccd1 _07719_/A sky130_fd_sc_hd__inv_2
XPHY_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _11836_/X _08685_/X _12702_/Q _08686_/X vssd1 vssd1 vccd1 vccd1 _12702_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ _12951_/Q vssd1 vssd1 vccd1 vccd1 _07649_/Y sky130_fd_sc_hd__inv_2
XPHY_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10660_ _08936_/A _08936_/B _09318_/A vssd1 vssd1 vccd1 vccd1 _10660_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09319_ _12370_/Q vssd1 vssd1 vccd1 vccd1 _09333_/A sky130_fd_sc_hd__inv_2
XFILLER_55_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10591_ _10525_/A _09390_/Y _09384_/Y vssd1 vssd1 vccd1 vccd1 _10591_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_103_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12330_ _12802_/CLK _12330_/D vssd1 vssd1 vccd1 vccd1 _12330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12261_ _12785_/Q _12858_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12261_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11212_ vssd1 vssd1 vccd1 vccd1 _11212_/HI _11212_/LO sky130_fd_sc_hd__conb_1
XFILLER_108_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12192_ _10790_/A _11145_/A _12193_/S vssd1 vssd1 vccd1 vccd1 _12192_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11143_ _10758_/A _10788_/A _13249_/Q _11111_/A _12116_/X vssd1 vssd1 vccd1 vccd1
+ _11143_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_132_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12664_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11074_ _10779_/X _11054_/X _06389_/X _11055_/X _11060_/X vssd1 vssd1 vccd1 vccd1
+ _11074_/X sky130_fd_sc_hd__a221o_1
Xinput120 la_data_in[58] vssd1 vssd1 vccd1 vccd1 input120/X sky130_fd_sc_hd__buf_1
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput131 la_data_in[68] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_hd__buf_1
XFILLER_49_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput142 la_data_in[78] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_hd__buf_1
X_10025_ _10168_/A vssd1 vssd1 vccd1 vccd1 _10025_/X sky130_fd_sc_hd__clkbuf_2
Xinput153 la_data_in[88] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_hd__buf_1
XFILLER_37_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput164 la_data_in[98] vssd1 vssd1 vccd1 vccd1 input164/X sky130_fd_sc_hd__buf_1
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput175 la_oenb[107] vssd1 vssd1 vccd1 vccd1 input175/X sky130_fd_sc_hd__buf_1
XFILLER_49_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput186 la_oenb[117] vssd1 vssd1 vccd1 vccd1 input186/X sky130_fd_sc_hd__buf_1
Xinput197 la_oenb[127] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__buf_1
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11976_ _10128_/Y _12792_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11976_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10927_ _10947_/A _10926_/X _10947_/A _10926_/X vssd1 vssd1 vccd1 vccd1 _12342_/D
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_177_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10858_ _10858_/A vssd1 vssd1 vccd1 vccd1 _10864_/C sky130_fd_sc_hd__inv_2
XFILLER_198_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _10736_/X _10788_/X _13252_/Q _10732_/X _10733_/X vssd1 vssd1 vccd1 vccd1
+ _10789_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12528_ _12535_/CLK _12528_/D vssd1 vssd1 vccd1 vccd1 _12528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12459_ _12978_/CLK _12459_/D vssd1 vssd1 vccd1 vccd1 _12459_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput605 _12291_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_67_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06951_ _06829_/X _09576_/B _06459_/X _06950_/X vssd1 vssd1 vccd1 vccd1 _13181_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09670_ _09668_/A _09668_/B _09669_/Y vssd1 vssd1 vccd1 vccd1 _09671_/B sky130_fd_sc_hd__a21o_1
X_06882_ _06890_/A _06890_/B vssd1 vssd1 vccd1 vccd1 _06883_/B sky130_fd_sc_hd__and2_1
XFILLER_95_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08621_ _08623_/A vssd1 vssd1 vccd1 vccd1 _08621_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08552_ _08550_/X _08552_/B vssd1 vssd1 vccd1 vccd1 _08552_/X sky130_fd_sc_hd__and2b_1
XFILLER_78_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07503_ _09184_/B vssd1 vssd1 vccd1 vccd1 _09227_/B sky130_fd_sc_hd__inv_2
XFILLER_51_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08483_ _13044_/Q _07823_/Y _13067_/Q _07824_/Y vssd1 vssd1 vccd1 vccd1 _08483_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07434_ _11474_/X _07429_/X _13033_/Q _07430_/X vssd1 vssd1 vccd1 vccd1 _13033_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07365_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07365_/X sky130_fd_sc_hd__clkbuf_1
X_09104_ _12532_/Q _09099_/X _09179_/D _09100_/X vssd1 vssd1 vccd1 vccd1 _12532_/D
+ sky130_fd_sc_hd__a22o_1
X_06316_ _06316_/A vssd1 vssd1 vccd1 vccd1 _06316_/X sky130_fd_sc_hd__clkbuf_4
X_07296_ _09186_/A vssd1 vssd1 vccd1 vccd1 _07296_/X sky130_fd_sc_hd__buf_2
XFILLER_175_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09035_ _09284_/A _09035_/B vssd1 vssd1 vccd1 vccd1 _09036_/B sky130_fd_sc_hd__or2_1
X_06247_ _06281_/A vssd1 vssd1 vccd1 vccd1 _06247_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06178_ _06174_/Y _06130_/B _06320_/A _06177_/X vssd1 vssd1 vccd1 vccd1 _06179_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_117_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09937_ _12669_/Q vssd1 vssd1 vccd1 vccd1 _09937_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09868_ _09868_/A _09880_/A _09868_/C vssd1 vssd1 vccd1 vccd1 _09868_/X sky130_fd_sc_hd__or3_2
XFILLER_86_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08819_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08819_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09799_ _13223_/Q _13222_/Q _09826_/A vssd1 vssd1 vccd1 vccd1 _09800_/B sky130_fd_sc_hd__o21ai_2
XPHY_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _09924_/Y _12855_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11830_/X sky130_fd_sc_hd__mux2_1
XPHY_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _12104_/X _11760_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11761_/X sky130_fd_sc_hd__mux2_1
XPHY_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10712_ _13240_/Q _11111_/A _10693_/A _10788_/A _06448_/Y vssd1 vssd1 vccd1 vccd1
+ _11110_/A sky130_fd_sc_hd__o221a_1
XPHY_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11691_/X _11395_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12388_/D sky130_fd_sc_hd__mux2_1
XPHY_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10643_ _10643_/A vssd1 vssd1 vccd1 vccd1 _10643_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10574_ _10583_/A _10574_/B vssd1 vssd1 vccd1 vccd1 _10574_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12313_ _12987_/CLK _12313_/D vssd1 vssd1 vccd1 vccd1 _12313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12244_ _12243_/X _12642_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12244_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12175_ _11142_/X _11137_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _12175_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11126_ _10779_/A _11100_/X _13245_/Q _11107_/X _11108_/X vssd1 vssd1 vccd1 vccd1
+ _11126_/X sky130_fd_sc_hd__a221o_1
XFILLER_3_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11057_ _06383_/X _11045_/X _11032_/X _10767_/X _11034_/X vssd1 vssd1 vccd1 vccd1
+ _11057_/X sky130_fd_sc_hd__a32o_1
XFILLER_7_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10008_ _08756_/Y _10003_/X _06203_/Y _10000_/X _10001_/X vssd1 vssd1 vccd1 vccd1
+ _10008_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_37_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11959_ _06494_/A _11141_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _11959_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07150_ _07152_/A vssd1 vssd1 vccd1 vccd1 _07150_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06101_ _06099_/Y _06100_/Y _12725_/Q _12693_/Q vssd1 vssd1 vccd1 vccd1 _06102_/A
+ sky130_fd_sc_hd__o22a_1
X_07081_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07081_/X sky130_fd_sc_hd__buf_1
XFILLER_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput402 _10109_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__clkbuf_2
X_06032_ _12747_/Q vssd1 vssd1 vccd1 vccd1 _06032_/Y sky130_fd_sc_hd__inv_2
Xoutput413 _11195_/LO vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput424 _11205_/LO vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__clkbuf_2
Xoutput435 _11215_/LO vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput446 _11216_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput457 _11226_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput468 _11227_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput479 _11230_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07983_ _10528_/C vssd1 vssd1 vccd1 vccd1 _07983_/X sky130_fd_sc_hd__buf_2
XFILLER_86_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09722_ _06735_/Y _06739_/Y _09705_/Y _09706_/Y vssd1 vssd1 vccd1 vccd1 _09722_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06934_ _06938_/A _06938_/B vssd1 vssd1 vccd1 vccd1 _06935_/B sky130_fd_sc_hd__and2_1
XFILLER_67_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09653_ _09653_/A vssd1 vssd1 vccd1 vccd1 _09653_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06865_ _13190_/Q vssd1 vssd1 vccd1 vccd1 _06865_/Y sky130_fd_sc_hd__inv_2
X_08604_ _08606_/A vssd1 vssd1 vccd1 vccd1 _08604_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09584_ _12870_/Q vssd1 vssd1 vccd1 vccd1 _09584_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06796_ _13198_/Q vssd1 vssd1 vccd1 vccd1 _06796_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08535_ _08535_/A vssd1 vssd1 vccd1 vccd1 _10691_/B sky130_fd_sc_hd__clkbuf_4
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08466_ _13056_/Q _10357_/B _13070_/Q _10393_/A vssd1 vssd1 vccd1 vccd1 _08466_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07417_ _07462_/A vssd1 vssd1 vccd1 vccd1 _07428_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08397_ _08405_/A vssd1 vssd1 vccd1 vccd1 _08397_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07348_ _07360_/A vssd1 vssd1 vccd1 vccd1 _07348_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07279_ _11548_/X _07248_/A _13083_/Q _07249_/A vssd1 vssd1 vccd1 vccd1 _13083_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09018_ _09019_/A _09019_/B _11636_/X vssd1 vssd1 vccd1 vccd1 _12580_/D sky130_fd_sc_hd__and3_1
X_10290_ _10283_/Y _10038_/X _09629_/Y _10033_/X _10289_/X vssd1 vssd1 vccd1 vccd1
+ _10290_/X sky130_fd_sc_hd__o221a_1
XFILLER_191_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12931_ _12973_/CLK _12931_/D vssd1 vssd1 vccd1 vccd1 _12931_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_92_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12862_ _12864_/CLK _12862_/D _08059_/X vssd1 vssd1 vccd1 vccd1 _12862_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _09179_/D _11812_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11813_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12793_ _13146_/CLK _12793_/D _08383_/X vssd1 vssd1 vccd1 vccd1 _12793_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11744_ _09185_/D _11743_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11744_/X sky130_fd_sc_hd__mux2_1
XPHY_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _11385_/X _09185_/A _11675_/S vssd1 vssd1 vccd1 vccd1 _11675_/X sky130_fd_sc_hd__mux2_1
XPHY_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ _12321_/Q _08925_/B _10608_/A _12417_/Q vssd1 vssd1 vccd1 vccd1 _10627_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10557_ _11391_/X _10557_/B vssd1 vssd1 vccd1 vccd1 _10557_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13276_ _13276_/CLK _13276_/D _06235_/X vssd1 vssd1 vccd1 vccd1 _13276_/Q sky130_fd_sc_hd__dfrtp_1
X_10488_ input32/X vssd1 vssd1 vccd1 vccd1 _10488_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12227_ _06291_/Y _13159_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12227_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12158_ _10012_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12158_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11109_ _11033_/X _11100_/X _13243_/Q _11107_/X _11108_/X vssd1 vssd1 vccd1 vccd1
+ _11109_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13253_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12089_ _10704_/Y _06535_/A _12762_/Q vssd1 vssd1 vccd1 vccd1 _12089_/X sky130_fd_sc_hd__mux2_2
XFILLER_96_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06650_ _06650_/A vssd1 vssd1 vccd1 vccd1 _06650_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06581_ _13220_/Q vssd1 vssd1 vccd1 vccd1 _06581_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08320_ _08325_/A vssd1 vssd1 vccd1 vccd1 _08320_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08251_ _08251_/A vssd1 vssd1 vccd1 vccd1 _08251_/X sky130_fd_sc_hd__clkbuf_2
X_07202_ _07263_/A vssd1 vssd1 vccd1 vccd1 _07264_/A sky130_fd_sc_hd__inv_2
XFILLER_159_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08182_ _13120_/Q _10420_/A _08180_/Y _12818_/Q _08181_/X vssd1 vssd1 vccd1 vccd1
+ _08190_/B sky130_fd_sc_hd__o221a_1
XFILLER_158_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07133_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07133_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07064_ _07053_/X _07058_/X _06316_/X _13154_/Q _07059_/X vssd1 vssd1 vccd1 vccd1
+ _13154_/D sky130_fd_sc_hd__a32o_1
XFILLER_12_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06015_ _07750_/B vssd1 vssd1 vccd1 vccd1 _09282_/A sky130_fd_sc_hd__inv_2
XFILLER_160_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07966_ _07985_/A vssd1 vssd1 vccd1 vccd1 _07966_/X sky130_fd_sc_hd__clkbuf_1
X_09705_ _13206_/Q vssd1 vssd1 vccd1 vccd1 _09705_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06917_ _06917_/A vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__clkbuf_2
X_07897_ _07903_/A vssd1 vssd1 vccd1 vccd1 _07897_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09636_ _13193_/Q _13192_/Q _09635_/Y _06844_/Y vssd1 vssd1 vccd1 vccd1 _09638_/A
+ sky130_fd_sc_hd__o22a_1
X_06848_ _12015_/X _06846_/B _06846_/X vssd1 vssd1 vccd1 vccd1 _06848_/X sky130_fd_sc_hd__a21bo_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09567_ _09568_/A _09568_/B vssd1 vssd1 vccd1 vccd1 _09567_/X sky130_fd_sc_hd__or2_1
X_06779_ _06719_/X _06774_/X _06778_/Y _06480_/X _13200_/Q vssd1 vssd1 vccd1 vccd1
+ _13200_/D sky130_fd_sc_hd__a32o_1
XFILLER_128_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08518_ _08518_/A vssd1 vssd1 vccd1 vccd1 _08518_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_196_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ _13170_/Q vssd1 vssd1 vccd1 vccd1 _09500_/A sky130_fd_sc_hd__inv_2
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08449_ _08445_/Y _07800_/X _08446_/Y _10388_/A _08448_/X vssd1 vssd1 vccd1 vccd1
+ _08457_/B sky130_fd_sc_hd__a221o_1
XPHY_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11460_ _12903_/Q _09243_/C _11469_/S vssd1 vssd1 vccd1 vccd1 _11460_/X sky130_fd_sc_hd__mux2_1
XPHY_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10411_ _10411_/A vssd1 vssd1 vccd1 vccd1 _10474_/A sky130_fd_sc_hd__buf_4
XFILLER_183_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11391_ _09333_/A _10555_/X _12321_/Q vssd1 vssd1 vccd1 vccd1 _11391_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13130_ _12168_/X _13130_/D _07152_/X vssd1 vssd1 vccd1 vccd1 _13130_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10342_ _10342_/A _10342_/B _10342_/C vssd1 vssd1 vccd1 vccd1 _10346_/C sky130_fd_sc_hd__or3_4
XFILLER_87_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13061_ _12165_/X _13061_/D _07352_/X vssd1 vssd1 vccd1 vccd1 _13061_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10273_ _10266_/Y _10038_/X _10267_/Y _10033_/X _10272_/X vssd1 vssd1 vccd1 vccd1
+ _10273_/X sky130_fd_sc_hd__o221a_1
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12012_ _11096_/X _11091_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _12012_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12576_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_94_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12914_ _12166_/X _12914_/D _07915_/X vssd1 vssd1 vccd1 vccd1 _12914_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12845_ _12864_/CLK _12845_/D _08103_/X vssd1 vssd1 vccd1 vccd1 _12845_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_73_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12776_ _12779_/CLK _12776_/D _08429_/X vssd1 vssd1 vccd1 vccd1 _12776_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11922_/X _12486_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11727_/X sky130_fd_sc_hd__mux2_1
XPHY_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _10557_/Y _10556_/Y _11704_/S vssd1 vssd1 vccd1 vccd1 _12370_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10609_ _10611_/A _10611_/B _10619_/A _09399_/Y vssd1 vssd1 vccd1 vccd1 _11888_/S
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11589_ _10432_/X _09243_/C _11592_/S vssd1 vssd1 vccd1 vccd1 _11589_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_1_wb_clk_i clkbuf_2_2_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13259_ _13260_/CLK _13259_/D _06329_/X vssd1 vssd1 vccd1 vccd1 _13259_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07820_ _13017_/Q vssd1 vssd1 vccd1 vccd1 _07820_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07751_ _08556_/B _12941_/Q _07751_/S vssd1 vssd1 vccd1 vccd1 _12941_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06702_ _06700_/X _06701_/X _06700_/X _06701_/X vssd1 vssd1 vccd1 vccd1 _06702_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07682_ _07682_/A vssd1 vssd1 vccd1 vccd1 _07682_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09421_ _12460_/Q _09411_/Y _12451_/Q _10525_/A _09420_/X vssd1 vssd1 vccd1 vccd1
+ _09421_/X sky130_fd_sc_hd__o221a_1
X_06633_ _12756_/Q _12757_/Q vssd1 vssd1 vccd1 vccd1 _06634_/A sky130_fd_sc_hd__and2_1
XFILLER_198_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _09349_/Y _12413_/Q _12456_/Q _09350_/Y _09351_/X vssd1 vssd1 vccd1 vccd1
+ _09353_/D sky130_fd_sc_hd__o221a_1
XFILLER_52_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06564_ _12174_/X _12173_/X _06562_/X vssd1 vssd1 vccd1 vccd1 _06564_/X sky130_fd_sc_hd__a21bo_1
XFILLER_33_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08303_ _12826_/Q _11601_/X _08307_/S vssd1 vssd1 vccd1 vccd1 _12826_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09283_ _09283_/A _09283_/B _09036_/B vssd1 vssd1 vccd1 vccd1 _12299_/D sky130_fd_sc_hd__or3b_2
X_06495_ _12042_/X vssd1 vssd1 vccd1 vccd1 _06495_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08234_ _08226_/Y _10405_/A _13107_/Q _08154_/Y vssd1 vssd1 vccd1 vccd1 _08237_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_178_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08165_ _13119_/Q vssd1 vssd1 vccd1 vccd1 _08165_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07116_ _07161_/A vssd1 vssd1 vccd1 vccd1 _07116_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_180_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08096_ _08098_/A vssd1 vssd1 vccd1 vccd1 _08096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07047_ _07037_/X _07040_/X _06283_/Y _13160_/Q _07042_/X vssd1 vssd1 vccd1 vccd1
+ _13160_/D sky130_fd_sc_hd__a32o_1
XFILLER_162_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08998_ _12939_/Q _12937_/Q _12938_/Q _08997_/X _07522_/A vssd1 vssd1 vccd1 vccd1
+ _12596_/D sky130_fd_sc_hd__a221o_1
XFILLER_48_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07949_ _08038_/A vssd1 vssd1 vccd1 vccd1 _07961_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10960_ _10952_/Y _10953_/Y _10977_/D _10977_/A vssd1 vssd1 vccd1 vccd1 _10960_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_141_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09619_ _13191_/Q _09618_/A _09617_/Y _09618_/Y vssd1 vssd1 vccd1 vccd1 _09620_/B
+ sky130_fd_sc_hd__a22o_1
X_10891_ _10873_/Y _10889_/X _10890_/Y _12524_/Q _12336_/Q vssd1 vssd1 vccd1 vccd1
+ _10891_/X sky130_fd_sc_hd__o32a_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12630_ _13170_/CLK _12630_/D _08895_/X vssd1 vssd1 vccd1 vccd1 _12630_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_157_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12344_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _12570_/CLK _12561_/D vssd1 vssd1 vccd1 vccd1 _12561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11512_ _10398_/X _10793_/B _11513_/S vssd1 vssd1 vccd1 vccd1 _11512_/X sky130_fd_sc_hd__mux2_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12492_ _12492_/CLK _12492_/D vssd1 vssd1 vccd1 vccd1 _12492_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11443_ _12918_/Q _10792_/A _11443_/S vssd1 vssd1 vccd1 vccd1 _11443_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11374_ _11373_/X _12427_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _11374_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ _12167_/X _13113_/D _07194_/X vssd1 vssd1 vccd1 vccd1 _13113_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10325_ _10325_/A _10326_/B _10387_/A vssd1 vssd1 vccd1 vccd1 _10325_/Y sky130_fd_sc_hd__nor3_2
XFILLER_153_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13044_ _12165_/X _13044_/D _07396_/X vssd1 vssd1 vccd1 vccd1 _13044_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10256_ _10254_/Y _10166_/X _10255_/Y _10168_/X vssd1 vssd1 vccd1 vccd1 _10256_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10187_ _10182_/Y _10163_/X _10183_/Y _10165_/X _10186_/X vssd1 vssd1 vccd1 vccd1
+ _10187_/X sky130_fd_sc_hd__o221a_1
XFILLER_94_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12828_ _12169_/X _12828_/D _08296_/X vssd1 vssd1 vccd1 vccd1 _12828_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12986_/CLK _12759_/D _08524_/X vssd1 vssd1 vccd1 vccd1 _12759_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06280_ _06280_/A vssd1 vssd1 vccd1 vccd1 _06280_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09970_ _10032_/A vssd1 vssd1 vccd1 vccd1 _09999_/A sky130_fd_sc_hd__buf_2
XFILLER_116_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08921_ _12420_/Q vssd1 vssd1 vccd1 vccd1 _08927_/A sky130_fd_sc_hd__inv_2
XFILLER_143_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08852_ _12615_/Q vssd1 vssd1 vccd1 vccd1 _08852_/X sky130_fd_sc_hd__buf_2
XFILLER_112_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07803_ _13016_/Q vssd1 vssd1 vccd1 vccd1 _07803_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08783_ _08789_/A vssd1 vssd1 vccd1 vccd1 _08783_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07734_ _07749_/A vssd1 vssd1 vccd1 vccd1 _07734_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07665_ _07665_/A _07665_/B _12956_/Q vssd1 vssd1 vccd1 vccd1 _07665_/X sky130_fd_sc_hd__and3_1
XFILLER_53_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09404_ _12409_/D vssd1 vssd1 vccd1 vccd1 _10603_/A sky130_fd_sc_hd__inv_2
X_06616_ _06616_/A vssd1 vssd1 vccd1 vccd1 _06620_/A sky130_fd_sc_hd__inv_2
XFILLER_197_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07596_ _09284_/A _09284_/B _12493_/Q _09288_/A _07595_/Y vssd1 vssd1 vccd1 vccd1
+ _12977_/D sky130_fd_sc_hd__o311a_1
XFILLER_111_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _12461_/Q vssd1 vssd1 vccd1 vccd1 _09335_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06547_ _12160_/X _11959_/X _06509_/Y _06510_/Y vssd1 vssd1 vccd1 vccd1 _06548_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_200_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09266_ _09434_/A _09434_/B vssd1 vssd1 vccd1 vccd1 _09266_/Y sky130_fd_sc_hd__nor2_1
X_06478_ _06522_/A vssd1 vssd1 vccd1 vccd1 _06478_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08217_ _13104_/Q vssd1 vssd1 vccd1 vccd1 _08217_/Y sky130_fd_sc_hd__inv_2
X_09197_ _12488_/Q _09190_/X _09180_/C _09192_/X vssd1 vssd1 vccd1 vccd1 _12488_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08148_ _13133_/Q _10454_/A _08147_/Y _12822_/Q vssd1 vssd1 vccd1 vccd1 _08151_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08079_ _08085_/A vssd1 vssd1 vccd1 vccd1 _08079_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10110_ _10109_/Y _10090_/X _08112_/Y _10047_/B vssd1 vssd1 vccd1 vccd1 _10110_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11090_ _10758_/X _11071_/X _06376_/X _11058_/X _11072_/X vssd1 vssd1 vccd1 vccd1
+ _11090_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput302 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__clkbuf_1
X_10041_ _10041_/A _10041_/B _10041_/C _10041_/D vssd1 vssd1 vccd1 vccd1 _10041_/Y
+ sky130_fd_sc_hd__nand4_2
Xinput313 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _07096_/A sky130_fd_sc_hd__clkbuf_1
Xinput324 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _09043_/A sky130_fd_sc_hd__buf_2
XFILLER_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput335 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 _07975_/A sky130_fd_sc_hd__buf_2
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput346 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 _10792_/A sky130_fd_sc_hd__buf_6
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput357 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 input357/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11992_ _11057_/X _11052_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _11992_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10943_ _10945_/D _10942_/X _10945_/D _10942_/X vssd1 vssd1 vccd1 vccd1 _12345_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10874_ _10873_/A _10873_/B _10873_/Y vssd1 vssd1 vccd1 vccd1 _10877_/A sky130_fd_sc_hd__a21oi_2
XFILLER_32_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12613_ _13162_/CLK _12614_/Q _08965_/X vssd1 vssd1 vccd1 vccd1 _12613_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12544_ _12547_/CLK _12544_/D vssd1 vssd1 vccd1 vccd1 _12544_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12475_ _12477_/CLK _12475_/D vssd1 vssd1 vccd1 vccd1 _12475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11426_ _12901_/Q _09183_/A _11433_/S vssd1 vssd1 vccd1 vccd1 _11426_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_54_wb_clk_i _12328_/CLK vssd1 vssd1 vccd1 vccd1 _12987_/CLK sky130_fd_sc_hd__clkbuf_16
X_11357_ _09331_/A _10549_/X _12321_/Q vssd1 vssd1 vccd1 vccd1 _11357_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10308_ _13096_/Q _10276_/X _13128_/Q _10277_/X vssd1 vssd1 vccd1 vccd1 _10308_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11288_ vssd1 vssd1 vccd1 vccd1 _11288_/HI _11288_/LO sky130_fd_sc_hd__conb_1
XFILLER_193_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13027_ _12164_/X _13027_/D _07448_/X vssd1 vssd1 vccd1 vccd1 _13027_/Q sky130_fd_sc_hd__dfrtp_4
X_10239_ _12648_/Q vssd1 vssd1 vccd1 vccd1 _10239_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07450_ _07458_/A vssd1 vssd1 vccd1 vccd1 _07450_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06401_ _06382_/X _12210_/X _06396_/X _06400_/X vssd1 vssd1 vccd1 vccd1 _13242_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_195_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07381_ _07391_/A vssd1 vssd1 vccd1 vccd1 _07381_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09120_ _12520_/Q _09115_/X _07993_/X _09116_/X vssd1 vssd1 vccd1 vccd1 _12520_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06332_ _06332_/A vssd1 vssd1 vccd1 vccd1 _06332_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_175_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09051_ _09051_/A _12154_/X vssd1 vssd1 vccd1 vccd1 _12565_/D sky130_fd_sc_hd__nor2b_1
X_06263_ _13271_/Q vssd1 vssd1 vccd1 vccd1 _06263_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08002_ _08004_/A vssd1 vssd1 vccd1 vccd1 _08002_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06194_ _06214_/A vssd1 vssd1 vccd1 vccd1 _06194_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09953_ _08774_/Y _09952_/X _06233_/X _09949_/X _09950_/X vssd1 vssd1 vccd1 vccd1
+ _09953_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_48_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08904_ _08898_/X _06327_/Y _08893_/X _12627_/Q vssd1 vssd1 vccd1 vccd1 _12627_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09884_ _09884_/A vssd1 vssd1 vccd1 vccd1 _09884_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08835_ _08814_/A _08781_/A _06351_/X _12654_/Q _08567_/A vssd1 vssd1 vccd1 vccd1
+ _12654_/D sky130_fd_sc_hd__a32o_1
XFILLER_58_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08766_ _08769_/A vssd1 vssd1 vccd1 vccd1 _08766_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ _07717_/A vssd1 vssd1 vccd1 vccd1 _07717_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _08699_/A vssd1 vssd1 vccd1 vccd1 _08697_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07648_ _07648_/A _07684_/B vssd1 vssd1 vccd1 vccd1 _07654_/B sky130_fd_sc_hd__or2_1
XPHY_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07579_ _12983_/Q _07574_/X _09185_/B _07575_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _12983_/D sky130_fd_sc_hd__o221a_1
XFILLER_55_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09318_ _09318_/A vssd1 vssd1 vccd1 vccd1 _12090_/S sky130_fd_sc_hd__inv_2
XFILLER_16_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10590_ _12403_/D _12404_/D _10525_/A _09390_/Y _11403_/S vssd1 vssd1 vccd1 vccd1
+ _10590_/X sky130_fd_sc_hd__o221a_1
XFILLER_51_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09249_ _12458_/Q _09251_/A _10528_/B _09083_/X vssd1 vssd1 vccd1 vccd1 _12458_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12260_ _12259_/X _12650_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12260_/X sky130_fd_sc_hd__mux2_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11211_ vssd1 vssd1 vccd1 vccd1 _11211_/HI _11211_/LO sky130_fd_sc_hd__conb_1
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12191_ _11139_/A _10782_/A _12193_/S vssd1 vssd1 vccd1 vccd1 _12191_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11142_ _10742_/A _11100_/A _13251_/Q _11107_/X _11108_/X vssd1 vssd1 vccd1 vccd1
+ _11142_/X sky130_fd_sc_hd__a221o_1
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11073_ _10767_/X _11071_/X _06383_/X _11058_/X _11072_/X vssd1 vssd1 vccd1 vccd1
+ _11073_/X sky130_fd_sc_hd__a221o_1
XFILLER_49_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput110 la_data_in[49] vssd1 vssd1 vccd1 vccd1 input110/X sky130_fd_sc_hd__buf_1
Xinput121 la_data_in[59] vssd1 vssd1 vccd1 vccd1 input121/X sky130_fd_sc_hd__buf_1
Xinput132 la_data_in[69] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_hd__buf_1
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10024_ _12638_/Q vssd1 vssd1 vccd1 vccd1 _10024_/Y sky130_fd_sc_hd__inv_2
Xinput143 la_data_in[79] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_hd__buf_1
XFILLER_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput154 la_data_in[89] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_hd__buf_1
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput165 la_data_in[99] vssd1 vssd1 vccd1 vccd1 input165/X sky130_fd_sc_hd__buf_1
Xinput176 la_oenb[108] vssd1 vssd1 vccd1 vccd1 input176/X sky130_fd_sc_hd__buf_1
Xinput187 la_oenb[118] vssd1 vssd1 vccd1 vccd1 input187/X sky130_fd_sc_hd__buf_1
XFILLER_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput198 la_oenb[12] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__buf_1
XFILLER_91_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_101_wb_clk_i _13235_/CLK vssd1 vssd1 vccd1 vccd1 _13236_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11975_ _10107_/Y _12791_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11975_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926_ _10895_/A _10944_/A _10947_/C vssd1 vssd1 vccd1 vccd1 _10926_/X sky130_fd_sc_hd__o21a_1
XFILLER_189_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10857_ _12520_/Q _12332_/Q _10851_/X _10852_/X vssd1 vssd1 vccd1 vccd1 _10859_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _10788_/A vssd1 vssd1 vccd1 vccd1 _10788_/X sky130_fd_sc_hd__clkbuf_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ _12529_/CLK _12527_/D vssd1 vssd1 vccd1 vccd1 _12527_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12458_ _12458_/CLK _12458_/D vssd1 vssd1 vccd1 vccd1 _12458_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput606 _12292_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__clkbuf_2
X_11409_ _12443_/Q _10659_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _11409_/X sky130_fd_sc_hd__mux2_1
X_12389_ _12413_/CLK _12389_/D vssd1 vssd1 vccd1 vccd1 _12411_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_181_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06950_ _06946_/X _06947_/X _06949_/X vssd1 vssd1 vccd1 vccd1 _06950_/X sky130_fd_sc_hd__o21a_1
XFILLER_141_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06881_ _12030_/X _06850_/X _12030_/X _06850_/X vssd1 vssd1 vccd1 vccd1 _06890_/B
+ sky130_fd_sc_hd__a2bb2oi_4
X_08620_ _11942_/X _08608_/X _12733_/Q _08610_/X vssd1 vssd1 vccd1 vccd1 _12733_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08551_ _12750_/Q _11963_/X _12610_/Q vssd1 vssd1 vccd1 vccd1 _08552_/B sky130_fd_sc_hd__o21ai_1
XFILLER_36_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07502_ _07609_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _13008_/D sky130_fd_sc_hd__nor2_1
XFILLER_78_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08482_ _08476_/X _08482_/B _08482_/C _08482_/D vssd1 vssd1 vccd1 vccd1 _08494_/C
+ sky130_fd_sc_hd__and4b_1
X_07433_ _07443_/A vssd1 vssd1 vccd1 vccd1 _07433_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07364_ _11433_/X _07353_/X _13057_/Q _07354_/X vssd1 vssd1 vccd1 vccd1 _13057_/D
+ sky130_fd_sc_hd__a22o_1
X_09103_ _12533_/Q _09099_/X _09179_/C _09100_/X vssd1 vssd1 vccd1 vccd1 _12533_/D
+ sky130_fd_sc_hd__a22o_1
X_06315_ _06129_/A _06103_/B _06130_/C _06102_/A vssd1 vssd1 vccd1 vccd1 _06316_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_175_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07295_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07295_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09034_ _13007_/Q _09284_/B _09276_/B vssd1 vssd1 vccd1 vccd1 _09035_/B sky130_fd_sc_hd__o21a_1
XFILLER_175_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06246_ _13274_/Q vssd1 vssd1 vccd1 vccd1 _06246_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06177_ _06098_/A _06102_/A _06176_/Y _06094_/X vssd1 vssd1 vccd1 vccd1 _06177_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_105_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09936_ _09934_/Y _09922_/X _06278_/A _09915_/X _09935_/X vssd1 vssd1 vccd1 vccd1
+ _09936_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09867_ _09828_/X _09868_/A _09839_/X vssd1 vssd1 vccd1 vccd1 _09867_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08818_ _08814_/X _08817_/X _06311_/Y _12662_/Q _08811_/X vssd1 vssd1 vccd1 vccd1
+ _12662_/D sky130_fd_sc_hd__a32o_1
XFILLER_93_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09798_ _09798_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__or2_2
XPHY_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _08748_/Y _08565_/X _06192_/X _08742_/X vssd1 vssd1 vccd1 vccd1 _12683_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_199_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _09185_/B _11759_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11760_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _10711_/A vssd1 vssd1 vccd1 vccd1 _10788_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _11395_/X _10528_/B _11691_/S vssd1 vssd1 vccd1 vccd1 _11691_/X sky130_fd_sc_hd__mux2_1
XPHY_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _11904_/X _10649_/B vssd1 vssd1 vccd1 vccd1 _10642_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10573_ _12399_/D _11390_/S _10520_/C _10564_/A vssd1 vssd1 vccd1 vccd1 _10574_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12312_ _12550_/CLK _12312_/D vssd1 vssd1 vccd1 vccd1 _12312_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_154_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12243_ _12776_/Q _12849_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12243_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12174_ _11136_/X _11132_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12174_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ _10767_/X _10759_/A _13247_/Q _11086_/X _11087_/X vssd1 vssd1 vccd1 vccd1
+ _11125_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11056_ _10699_/X _11054_/X _06400_/X _11055_/X _10747_/X vssd1 vssd1 vccd1 vccd1
+ _11056_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10007_ _08759_/Y _10003_/X _06207_/Y _10000_/X _10001_/X vssd1 vssd1 vccd1 vccd1
+ _10007_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11958_ _09886_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11958_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10909_ _12527_/Q _12339_/Q _10900_/Y _10904_/A vssd1 vssd1 vccd1 vccd1 _10909_/X
+ sky130_fd_sc_hd__o22a_1
X_11889_ _10625_/Y _12416_/D _11889_/S vssd1 vssd1 vccd1 vccd1 _11889_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06100_ _12693_/Q vssd1 vssd1 vccd1 vccd1 _06100_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07080_ _07154_/A vssd1 vssd1 vccd1 vccd1 _07122_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06031_ _12748_/Q _12716_/Q _12748_/Q _12716_/Q vssd1 vssd1 vccd1 vccd1 _06035_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_201_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput403 _12965_/Q vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_201_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput414 _11196_/LO vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput425 _11206_/LO vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput436 _11185_/LO vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput447 _11316_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput458 _11326_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput469 _11336_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__clkbuf_2
XFILLER_102_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07982_ _07985_/A vssd1 vssd1 vccd1 vccd1 _07982_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09721_ _13210_/Q vssd1 vssd1 vccd1 vccd1 _09721_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06933_ _12028_/X _06902_/X _12028_/X _06902_/X vssd1 vssd1 vccd1 vccd1 _06938_/B
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_80_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09652_ _13197_/Q vssd1 vssd1 vccd1 vccd1 _09652_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06864_ _06864_/A _06864_/B vssd1 vssd1 vccd1 vccd1 _06864_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08603_ _11948_/X _08592_/X _12739_/Q _08593_/X vssd1 vssd1 vccd1 vccd1 _12739_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09583_ _09582_/A _09582_/B _09701_/A vssd1 vssd1 vccd1 vccd1 _09583_/Y sky130_fd_sc_hd__o21ai_1
X_06795_ _06806_/A vssd1 vssd1 vccd1 vccd1 _06795_/X sky130_fd_sc_hd__clkbuf_1
X_08534_ _12755_/Q vssd1 vssd1 vccd1 vccd1 _08535_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08465_ _13061_/Q _10367_/A _08464_/Y _12911_/Q vssd1 vssd1 vccd1 vccd1 _08467_/C
+ sky130_fd_sc_hd__a22o_1
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07416_ _11481_/X _07412_/X _13040_/Q _07415_/X vssd1 vssd1 vccd1 vccd1 _13040_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08396_ _12788_/Q _08374_/A _07313_/X _08375_/A vssd1 vssd1 vccd1 vccd1 _12788_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07347_ _07362_/A vssd1 vssd1 vccd1 vccd1 _07360_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07278_ _07280_/A vssd1 vssd1 vccd1 vccd1 _07278_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09017_ _09019_/A _09019_/B _11637_/X vssd1 vssd1 vccd1 vccd1 _12581_/D sky130_fd_sc_hd__and3_1
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06229_ _06227_/Y _06216_/X _06217_/X _06228_/X vssd1 vssd1 vccd1 vccd1 _13278_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_152_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09919_ _12886_/Q _09919_/B vssd1 vssd1 vccd1 vccd1 _09919_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12930_ _12937_/CLK _12930_/D vssd1 vssd1 vccd1 vccd1 _12930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12861_ _12864_/CLK _12861_/D _08061_/X vssd1 vssd1 vccd1 vccd1 _12861_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11812_ _12086_/X _12491_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11812_/X sky130_fd_sc_hd__mux2_1
XPHY_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _13146_/CLK _12792_/D _08385_/X vssd1 vssd1 vccd1 vccd1 _12792_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11372_/X _12470_/Q _12103_/S vssd1 vssd1 vccd1 vccd1 _11743_/X sky130_fd_sc_hd__mux2_1
XPHY_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _11673_/X _11387_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12379_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10625_ _10625_/A _11888_/X vssd1 vssd1 vccd1 vccd1 _10625_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10556_ _11391_/X vssd1 vssd1 vccd1 vccd1 _10556_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13275_ _13279_/CLK _13275_/D _06239_/X vssd1 vssd1 vccd1 vccd1 _13275_/Q sky130_fd_sc_hd__dfrtp_1
X_10487_ _12835_/Q _10486_/Y _08122_/Y _10486_/A _10459_/X vssd1 vssd1 vccd1 vccd1
+ _10487_/X sky130_fd_sc_hd__o221a_1
XFILLER_154_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12226_ _12225_/X _12633_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12226_/X sky130_fd_sc_hd__mux2_2
XFILLER_194_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12157_ _10011_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12157_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ _12132_/X vssd1 vssd1 vccd1 vccd1 _11108_/X sky130_fd_sc_hd__clkbuf_2
X_12088_ _06634_/A _10701_/Y _12758_/Q vssd1 vssd1 vccd1 vccd1 _12186_/S sky130_fd_sc_hd__mux2_8
XFILLER_110_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11039_ _10696_/X _11037_/X _06404_/X _07020_/X _11038_/X vssd1 vssd1 vccd1 vccd1
+ _11039_/X sky130_fd_sc_hd__a221o_1
XFILLER_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06580_ _06580_/A vssd1 vssd1 vccd1 vccd1 _06580_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08250_ _08250_/A vssd1 vssd1 vccd1 vccd1 _11417_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07201_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07201_/X sky130_fd_sc_hd__clkbuf_2
X_08181_ _13131_/Q _12821_/Q _13131_/Q _12821_/Q vssd1 vssd1 vccd1 vccd1 _08181_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_146_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_wb_clk_i _12328_/CLK vssd1 vssd1 vccd1 vccd1 _12849_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07132_ _11540_/X _07130_/X _13139_/Q _07131_/X vssd1 vssd1 vccd1 vccd1 _13139_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07063_ _07063_/A vssd1 vssd1 vccd1 vccd1 _07063_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06014_ _12607_/Q _06017_/B _09259_/A vssd1 vssd1 vccd1 vccd1 _07750_/B sky130_fd_sc_hd__and3_1
XFILLER_160_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07965_ _10318_/A _11483_/X _07967_/S vssd1 vssd1 vccd1 vccd1 _12894_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09704_ _13205_/Q _13204_/Q _06735_/Y _06739_/Y vssd1 vssd1 vccd1 vccd1 _09706_/A
+ sky130_fd_sc_hd__o22a_1
X_06916_ _06916_/A vssd1 vssd1 vccd1 vccd1 _06916_/X sky130_fd_sc_hd__clkbuf_1
X_07896_ _10397_/A _11512_/X _07904_/S vssd1 vssd1 vccd1 vccd1 _12923_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09635_ _13193_/Q vssd1 vssd1 vccd1 vccd1 _09635_/Y sky130_fd_sc_hd__inv_2
X_06847_ _12025_/X _12021_/X _06846_/X vssd1 vssd1 vccd1 vccd1 _06847_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06778_ _06778_/A _06778_/B vssd1 vssd1 vccd1 vccd1 _06778_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09566_ _09566_/A _09566_/B vssd1 vssd1 vccd1 vccd1 _09568_/B sky130_fd_sc_hd__or2_1
XFILLER_43_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ _08504_/X _12250_/X _08514_/X _12762_/Q vssd1 vssd1 vccd1 vccd1 _12762_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09497_ _13167_/Q _13166_/Q _13168_/Q _09488_/X vssd1 vssd1 vccd1 vccd1 _09502_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_196_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08448_ _08446_/Y _10388_/A _08447_/Y _07804_/X vssd1 vssd1 vccd1 vccd1 _08448_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08379_ _08385_/A vssd1 vssd1 vccd1 vccd1 _08379_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10410_ _12805_/Q _12804_/Q _12806_/Q vssd1 vssd1 vccd1 vccd1 _10413_/B sky130_fd_sc_hd__and3_1
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _10576_/X _12400_/D _11390_/S vssd1 vssd1 vccd1 vccd1 _11390_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10341_ _10342_/B _10342_/C _10342_/A vssd1 vssd1 vccd1 vccd1 _10344_/A sky130_fd_sc_hd__o21a_1
XFILLER_192_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13060_ _12165_/X _13060_/D _07356_/X vssd1 vssd1 vccd1 vccd1 _13060_/Q sky130_fd_sc_hd__dfrtp_4
X_10272_ _10268_/Y _10163_/A _10269_/Y _10165_/A _10271_/X vssd1 vssd1 vccd1 vccd1
+ _10272_/X sky130_fd_sc_hd__o221a_1
XFILLER_180_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12011_ _11080_/X _11070_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _12011_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_wb_clk_i _13219_/CLK vssd1 vssd1 vccd1 vccd1 _13217_/CLK sky130_fd_sc_hd__clkbuf_16
X_12913_ _12166_/X _12913_/D _07917_/X vssd1 vssd1 vccd1 vccd1 _12913_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12844_ _12844_/CLK _12844_/D vssd1 vssd1 vccd1 vccd1 _12844_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12987_/CLK _12775_/D _08431_/X vssd1 vssd1 vccd1 vccd1 _12775_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11726_ _08556_/B _09259_/Y _12607_/Q vssd1 vssd1 vccd1 vccd1 _11726_/X sky130_fd_sc_hd__mux2_1
XPHY_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _10554_/Y _10553_/Y _11704_/S vssd1 vssd1 vccd1 vccd1 _12369_/D sky130_fd_sc_hd__mux2_1
XPHY_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10608_ _10608_/A _10608_/B _12371_/Q vssd1 vssd1 vccd1 vccd1 _11889_/S sky130_fd_sc_hd__or3b_4
XPHY_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11588_ _10431_/Y _09243_/D _11592_/S vssd1 vssd1 vccd1 vccd1 _11588_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10539_ _11360_/X vssd1 vssd1 vccd1 vccd1 _10539_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13258_ _13260_/CLK _13258_/D _06334_/X vssd1 vssd1 vccd1 vccd1 _13258_/Q sky130_fd_sc_hd__dfrtp_1
X_12209_ _06336_/Y _13150_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12209_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13189_ _13190_/CLK _13189_/D _06869_/X vssd1 vssd1 vccd1 vccd1 _13189_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_85_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07750_ _11726_/X _07750_/B vssd1 vssd1 vccd1 vccd1 _07751_/S sky130_fd_sc_hd__or2_1
XFILLER_38_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06701_ _11987_/X _11990_/X _11987_/X _11990_/X vssd1 vssd1 vccd1 vccd1 _06701_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07681_ _12307_/Q _07726_/B vssd1 vssd1 vccd1 vccd1 _07682_/A sky130_fd_sc_hd__nand2_1
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09420_ _12457_/Q _10603_/A _12456_/Q _10599_/B vssd1 vssd1 vccd1 vccd1 _09420_/X
+ sky130_fd_sc_hd__o22a_1
X_06632_ _11896_/X _06632_/B vssd1 vssd1 vccd1 vccd1 _06632_/X sky130_fd_sc_hd__or2_1
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09351_ _12453_/Q _12405_/Q _12453_/Q _12405_/Q vssd1 vssd1 vccd1 vccd1 _09351_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06563_ _12178_/X _12177_/X _06562_/X vssd1 vssd1 vccd1 vccd1 _06563_/X sky130_fd_sc_hd__o21a_1
XFILLER_166_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08302_ _08311_/A vssd1 vssd1 vccd1 vccd1 _08302_/X sky130_fd_sc_hd__clkbuf_1
X_09282_ _09282_/A _09282_/B vssd1 vssd1 vccd1 vccd1 _12607_/D sky130_fd_sc_hd__nand2_1
XFILLER_61_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06494_ _06494_/A vssd1 vssd1 vccd1 vccd1 _06494_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_opt_1_wb_clk_i clkbuf_opt_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_08233_ _13109_/Q _10477_/A _08206_/Y _12813_/Q vssd1 vssd1 vccd1 vccd1 _08233_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08164_ _12828_/Q vssd1 vssd1 vccd1 vccd1 _08164_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07115_ _07177_/A vssd1 vssd1 vccd1 vccd1 _07161_/A sky130_fd_sc_hd__buf_4
XFILLER_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08095_ _12849_/Q _08082_/X _07296_/X _08083_/X vssd1 vssd1 vccd1 vccd1 _12849_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07046_ _07046_/A vssd1 vssd1 vccd1 vccd1 _07046_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08997_ _12939_/Q _12937_/Q vssd1 vssd1 vccd1 vccd1 _08997_/X sky130_fd_sc_hd__or2_1
XFILLER_69_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07948_ _08657_/A vssd1 vssd1 vccd1 vccd1 _08038_/A sky130_fd_sc_hd__buf_2
XFILLER_29_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07879_ _07870_/X _07879_/B _07879_/C _07879_/D vssd1 vssd1 vccd1 vccd1 _07879_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09618_ _09618_/A vssd1 vssd1 vccd1 vccd1 _09618_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ _10890_/A _10890_/B _10890_/C vssd1 vssd1 vccd1 vccd1 _10890_/Y sky130_fd_sc_hd__nor3_1
XFILLER_71_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09549_ _13178_/Q vssd1 vssd1 vccd1 vccd1 _09550_/A sky130_fd_sc_hd__inv_2
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _12570_/CLK _12560_/D vssd1 vssd1 vccd1 vccd1 _12560_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11511_ _10396_/Y _10794_/A _11513_/S vssd1 vssd1 vccd1 vccd1 _11511_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12491_ _12492_/CLK _12491_/D vssd1 vssd1 vccd1 vccd1 _12491_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11442_ _12917_/Q _10792_/B _11443_/S vssd1 vssd1 vccd1 vccd1 _11442_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_126_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13283_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11373_ _10664_/X _12427_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10324_ _10324_/A vssd1 vssd1 vccd1 vccd1 _10387_/A sky130_fd_sc_hd__buf_6
X_13112_ _12167_/X _13112_/D _07206_/X vssd1 vssd1 vccd1 vccd1 _13112_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13043_ _12165_/X _13043_/D _07398_/X vssd1 vssd1 vccd1 vccd1 _13043_/Q sky130_fd_sc_hd__dfrtp_1
X_10255_ _12649_/Q vssd1 vssd1 vccd1 vccd1 _10255_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10186_ _10184_/Y _10166_/X _10185_/Y _10168_/X vssd1 vssd1 vccd1 vccd1 _10186_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12827_ _12169_/X _12827_/D _08300_/X vssd1 vssd1 vccd1 vccd1 _12827_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_201_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12986_/CLK _12758_/D _08526_/X vssd1 vssd1 vccd1 vccd1 _12758_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11709_ _10634_/Y _10635_/Y _11818_/S vssd1 vssd1 vccd1 vccd1 _11709_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12689_ _12719_/CLK _12689_/D _08729_/X vssd1 vssd1 vccd1 vccd1 _12689_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08920_ _12421_/Q vssd1 vssd1 vccd1 vccd1 _08928_/A sky130_fd_sc_hd__inv_2
XFILLER_131_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08851_ _08851_/A vssd1 vssd1 vccd1 vccd1 _08851_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07802_ _12919_/Q vssd1 vssd1 vccd1 vccd1 _10388_/A sky130_fd_sc_hd__buf_2
X_08782_ _08780_/Y _08781_/X _06243_/X _08764_/X vssd1 vssd1 vccd1 vccd1 _12674_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_133_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07733_ _06358_/X _07729_/X _07732_/X vssd1 vssd1 vccd1 vccd1 _12945_/D sky130_fd_sc_hd__o21a_1
XFILLER_77_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07664_ _07664_/A vssd1 vssd1 vccd1 vccd1 _07664_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09403_ _12413_/D vssd1 vssd1 vccd1 vccd1 _10619_/A sky130_fd_sc_hd__inv_2
X_06615_ _11894_/X _11892_/X _06609_/X _06610_/X _06614_/X vssd1 vssd1 vccd1 vccd1
+ _06616_/A sky130_fd_sc_hd__o32a_1
X_07595_ _09284_/A _09284_/B _08977_/B vssd1 vssd1 vccd1 vccd1 _07595_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09334_ _12450_/Q _12619_/Q vssd1 vssd1 vccd1 vccd1 _09334_/X sky130_fd_sc_hd__or2_4
X_06546_ _06546_/A vssd1 vssd1 vccd1 vccd1 _06552_/A sky130_fd_sc_hd__inv_2
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09265_ _11966_/X vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__inv_2
X_06477_ _06766_/A vssd1 vssd1 vccd1 vccd1 _06522_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08216_ _08213_/Y _12821_/Q _13099_/Q _10455_/A _08215_/X vssd1 vssd1 vccd1 vccd1
+ _08222_/B sky130_fd_sc_hd__a221o_1
X_09196_ _12489_/Q _09190_/X _09180_/B _09192_/X vssd1 vssd1 vccd1 vccd1 _12489_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ _13132_/Q vssd1 vssd1 vccd1 vccd1 _08147_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08078_ _12856_/Q _08066_/X _07990_/X _08068_/X vssd1 vssd1 vccd1 vccd1 _12856_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_161_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07029_ _07046_/A vssd1 vssd1 vccd1 vccd1 _07029_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10040_ _10031_/Y _10032_/X _09476_/Y _10033_/X _10039_/X vssd1 vssd1 vccd1 vccd1
+ _10041_/D sky130_fd_sc_hd__o221a_1
Xinput303 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 _07101_/B sky130_fd_sc_hd__clkbuf_1
Xinput314 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _07096_/D sky130_fd_sc_hd__clkbuf_1
Xinput325 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _09043_/B sky130_fd_sc_hd__buf_2
Xinput336 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 input336/X sky130_fd_sc_hd__buf_2
XFILLER_76_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput347 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 _10794_/D sky130_fd_sc_hd__buf_6
Xinput358 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 input358/X sky130_fd_sc_hd__buf_4
XFILLER_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11991_ _11129_/Y _11121_/X _12193_/S vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10942_ _10936_/Y _10937_/Y _10945_/C _10939_/Y vssd1 vssd1 vccd1 vccd1 _10942_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10873_ _10873_/A _10873_/B vssd1 vssd1 vccd1 vccd1 _10873_/Y sky130_fd_sc_hd__nor2_4
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12688_/CLK _12613_/Q _08966_/X vssd1 vssd1 vccd1 vccd1 _12612_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12543_ _13001_/CLK _12543_/D vssd1 vssd1 vccd1 vccd1 _12543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12474_ _12474_/CLK _12474_/D vssd1 vssd1 vccd1 vccd1 _12474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11425_ _12900_/Q input358/X _11433_/S vssd1 vssd1 vccd1 vccd1 _11425_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11356_ _09468_/X _12993_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _12320_/D sky130_fd_sc_hd__mux2_1
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10307_ _10312_/A _11925_/X vssd1 vssd1 vccd1 vccd1 _10307_/Y sky130_fd_sc_hd__nor2b_4
XFILLER_98_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11287_ vssd1 vssd1 vccd1 vccd1 _11287_/HI _11287_/LO sky130_fd_sc_hd__conb_1
XFILLER_112_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13026_ _12164_/X _13026_/D _07450_/X vssd1 vssd1 vccd1 vccd1 _13026_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_94_wb_clk_i _12726_/CLK vssd1 vssd1 vccd1 vccd1 _13162_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10238_ _12632_/Q vssd1 vssd1 vccd1 vccd1 _10238_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12477_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10169_ _09535_/Y _10166_/X _10167_/Y _10168_/X vssd1 vssd1 vccd1 vccd1 _10169_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_66_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06400_ _13242_/Q vssd1 vssd1 vccd1 vccd1 _06400_/X sky130_fd_sc_hd__buf_2
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07380_ _11427_/X _07368_/X _13051_/Q _07369_/X vssd1 vssd1 vccd1 vccd1 _13051_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06331_ _06125_/A _06330_/X _06125_/A _06330_/X vssd1 vssd1 vccd1 vccd1 _06332_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_188_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09050_ _09051_/A _12155_/X vssd1 vssd1 vccd1 vccd1 _12566_/D sky130_fd_sc_hd__nor2b_1
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06262_ _06280_/A vssd1 vssd1 vccd1 vccd1 _06262_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08001_ _12885_/Q _07996_/X _07287_/X _07998_/X vssd1 vssd1 vccd1 vccd1 _12885_/D
+ sky130_fd_sc_hd__a22o_1
X_06193_ _06191_/Y _06022_/X _06163_/X _06192_/X vssd1 vssd1 vccd1 vccd1 _13284_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_144_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09952_ _09952_/A vssd1 vssd1 vccd1 vccd1 _09952_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08903_ _08912_/A vssd1 vssd1 vccd1 vccd1 _08903_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_131_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09883_ _09851_/B _09881_/B _09808_/B _09881_/X _09882_/X vssd1 vssd1 vccd1 vccd1
+ _09884_/A sky130_fd_sc_hd__o311a_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08834_ _08836_/A vssd1 vssd1 vccd1 vccd1 _08834_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08765_ _08763_/Y _08760_/X _06218_/X _08764_/X vssd1 vssd1 vccd1 vccd1 _12679_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_54_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _12952_/Q _07707_/X _12951_/Q _07705_/X _07714_/X vssd1 vssd1 vccd1 vccd1
+ _12952_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _11837_/X _08685_/X _12703_/Q _08686_/X vssd1 vssd1 vccd1 vccd1 _12703_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07647_ _12959_/Q _07652_/A _12958_/Q vssd1 vssd1 vccd1 vccd1 _07684_/B sky130_fd_sc_hd__nor3b_4
XPHY_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07578_ _12984_/Q _07574_/X _07536_/X _07575_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _12984_/D sky130_fd_sc_hd__o221a_1
XFILLER_16_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09317_ _12444_/Q _12443_/Q vssd1 vssd1 vccd1 vccd1 _09317_/X sky130_fd_sc_hd__or2_1
XFILLER_139_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06529_ _13225_/Q vssd1 vssd1 vccd1 vccd1 _06529_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09248_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09251_/A sky130_fd_sc_hd__inv_2
XFILLER_166_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09179_ _09179_/A _09179_/B _09179_/C _09179_/D vssd1 vssd1 vccd1 vccd1 _09187_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_147_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11210_ vssd1 vssd1 vccd1 vccd1 _11210_/HI _11210_/LO sky130_fd_sc_hd__conb_1
X_12190_ _10781_/A _10719_/X _12193_/S vssd1 vssd1 vccd1 vccd1 _12190_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11141_ _10730_/A _10759_/A _13253_/Q _11086_/A _12195_/X vssd1 vssd1 vccd1 vccd1
+ _11141_/X sky130_fd_sc_hd__a221o_1
XFILLER_150_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11072_ _12087_/X vssd1 vssd1 vccd1 vccd1 _11072_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput100 la_data_in[3] vssd1 vssd1 vccd1 vccd1 input100/X sky130_fd_sc_hd__buf_1
XFILLER_131_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput111 la_data_in[4] vssd1 vssd1 vccd1 vccd1 input111/X sky130_fd_sc_hd__buf_1
XFILLER_88_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput122 la_data_in[5] vssd1 vssd1 vccd1 vccd1 input122/X sky130_fd_sc_hd__buf_1
XFILLER_1_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10023_ _10166_/A vssd1 vssd1 vccd1 vccd1 _10023_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput133 la_data_in[6] vssd1 vssd1 vccd1 vccd1 input133/X sky130_fd_sc_hd__buf_1
Xinput144 la_data_in[7] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_hd__buf_1
Xinput155 la_data_in[8] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__buf_1
Xinput166 la_data_in[9] vssd1 vssd1 vccd1 vccd1 input166/X sky130_fd_sc_hd__buf_1
Xinput177 la_oenb[109] vssd1 vssd1 vccd1 vccd1 input177/X sky130_fd_sc_hd__buf_1
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput188 la_oenb[119] vssd1 vssd1 vccd1 vccd1 input188/X sky130_fd_sc_hd__buf_1
Xinput199 la_oenb[13] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__buf_1
XFILLER_5_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11974_ _10088_/Y _12790_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11974_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10925_ _10911_/Y _10912_/Y _10922_/X _10924_/Y vssd1 vssd1 vccd1 vccd1 _10947_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_141_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12942_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10856_ _12521_/Q _12333_/Q _10854_/Y _10855_/Y vssd1 vssd1 vccd1 vccd1 _10858_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10787_/A vssd1 vssd1 vccd1 vccd1 _10787_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _12529_/CLK _12526_/D vssd1 vssd1 vccd1 vccd1 _12526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12457_ _12547_/CLK _12457_/D vssd1 vssd1 vccd1 vccd1 _12457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11408_ _11049_/Y _10750_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _11408_/X sky130_fd_sc_hd__mux2_1
X_12388_ _12619_/CLK _12388_/D vssd1 vssd1 vccd1 vccd1 _12410_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11339_ vssd1 vssd1 vccd1 vccd1 _11339_/HI _11339_/LO sky130_fd_sc_hd__conb_1
XFILLER_67_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13009_ _12164_/X _13009_/D _07492_/X vssd1 vssd1 vccd1 vccd1 _13009_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06880_ _06873_/X _06877_/X _06883_/A vssd1 vssd1 vccd1 vccd1 _06890_/A sky130_fd_sc_hd__a21oi_4
XFILLER_95_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08550_ _12609_/Q _12608_/Q _12751_/Q _11963_/X vssd1 vssd1 vccd1 vccd1 _08550_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07501_ _09228_/A _07497_/Y _07522_/B _09279_/C _11982_/X vssd1 vssd1 vccd1 vccd1
+ _07502_/B sky130_fd_sc_hd__o32a_1
XFILLER_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08481_ _08447_/Y _07804_/X _13073_/Q _07809_/Y _08480_/Y vssd1 vssd1 vccd1 vccd1
+ _08482_/D sky130_fd_sc_hd__o221a_1
XFILLER_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07432_ _07462_/A vssd1 vssd1 vccd1 vccd1 _07443_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_189_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07363_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07363_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09102_ _12534_/Q _09099_/X _10792_/B _09100_/X vssd1 vssd1 vccd1 vccd1 _12534_/D
+ sky130_fd_sc_hd__a22o_1
X_06314_ _06314_/A vssd1 vssd1 vccd1 vccd1 _06314_/X sky130_fd_sc_hd__clkbuf_2
X_07294_ _07293_/X _07285_/X _07106_/X vssd1 vssd1 vccd1 vccd1 _13079_/D sky130_fd_sc_hd__o21a_1
X_09033_ _12300_/Q vssd1 vssd1 vccd1 vccd1 _09276_/B sky130_fd_sc_hd__inv_2
X_06245_ _06245_/A vssd1 vssd1 vccd1 vccd1 _06245_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06176_ _06176_/A vssd1 vssd1 vccd1 vccd1 _06176_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09935_ _12891_/Q _09935_/B vssd1 vssd1 vccd1 vccd1 _09935_/X sky130_fd_sc_hd__or2_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09866_ _09866_/A _09866_/B vssd1 vssd1 vccd1 vccd1 _09880_/A sky130_fd_sc_hd__or2_1
XFILLER_58_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08817_ _08817_/A vssd1 vssd1 vccd1 vccd1 _08817_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09797_ _06581_/Y _09787_/X _06577_/Y _09788_/X vssd1 vssd1 vccd1 vccd1 _09800_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _12683_/Q vssd1 vssd1 vccd1 vccd1 _08748_/Y sky130_fd_sc_hd__inv_2
XPHY_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _11844_/X _08670_/X _12710_/Q _08671_/X vssd1 vssd1 vccd1 vccd1 _12710_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _12767_/Q _12766_/Q vssd1 vssd1 vccd1 vccd1 _10710_/Y sky130_fd_sc_hd__nor2_2
XPHY_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11689_/X _11398_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12387_/D sky130_fd_sc_hd__mux2_1
XPHY_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10641_ _11904_/X vssd1 vssd1 vccd1 vccd1 _10641_/Y sky130_fd_sc_hd__inv_2
XPHY_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10572_ _10579_/A _10571_/Y _09415_/Y _10526_/A vssd1 vssd1 vccd1 vccd1 _10583_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_167_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12311_ _12951_/CLK _12311_/D vssd1 vssd1 vccd1 vccd1 _12311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12242_ _12241_/X _12641_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12242_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ _11135_/Y _11131_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _12173_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11124_ _10758_/X _11075_/A _06376_/X _11083_/X _11084_/X vssd1 vssd1 vccd1 vccd1
+ _11124_/X sky130_fd_sc_hd__a221o_1
XFILLER_122_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11055_ _11055_/A vssd1 vssd1 vccd1 vccd1 _11055_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10006_ _08763_/Y _10003_/X _06215_/Y _10000_/X _10001_/X vssd1 vssd1 vccd1 vccd1
+ _10006_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_77_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11957_ _09878_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11957_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10908_ _12528_/Q _12340_/Q _10906_/Y _10907_/Y vssd1 vssd1 vccd1 vccd1 _10908_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_72_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11888_ _10624_/X _10610_/B _11888_/S vssd1 vssd1 vccd1 vccd1 _11888_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10839_ _10837_/Y _10838_/Y _12518_/Q _12330_/Q vssd1 vssd1 vccd1 vccd1 _10864_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12509_ _12509_/CLK _12509_/D vssd1 vssd1 vccd1 vccd1 _12509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06030_ _06030_/A _06029_/Y vssd1 vssd1 vccd1 vccd1 _06185_/A sky130_fd_sc_hd__or2b_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput404 _11150_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__clkbuf_2
Xoutput415 _11197_/LO vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput426 _11207_/LO vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput437 _11346_/X vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput448 _11317_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput459 _11327_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07981_ _12891_/Q _07974_/X _07980_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _12891_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09720_ _09701_/X _09718_/X _09719_/Y _09682_/X vssd1 vssd1 vccd1 vccd1 _09720_/X
+ sky130_fd_sc_hd__a31o_1
X_06932_ _06925_/X _06929_/X _06935_/A vssd1 vssd1 vccd1 vccd1 _06938_/A sky130_fd_sc_hd__a21oi_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09651_ _13196_/Q _13195_/Q _06822_/Y _06830_/Y vssd1 vssd1 vccd1 vccd1 _09653_/A
+ sky130_fd_sc_hd__o22a_1
X_06863_ _06863_/A vssd1 vssd1 vccd1 vccd1 _06863_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08602_ _08606_/A vssd1 vssd1 vccd1 vccd1 _08602_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09582_ _09582_/A _09582_/B vssd1 vssd1 vccd1 vccd1 _09592_/B sky130_fd_sc_hd__and2_1
X_06794_ _06794_/A vssd1 vssd1 vccd1 vccd1 _13199_/D sky130_fd_sc_hd__inv_2
XFILLER_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08533_ _08533_/A vssd1 vssd1 vccd1 vccd1 _08533_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08464_ _13060_/Q vssd1 vssd1 vccd1 vccd1 _08464_/Y sky130_fd_sc_hd__inv_2
XPHY_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07415_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07415_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ _08405_/A vssd1 vssd1 vccd1 vccd1 _08395_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07346_ _11440_/X _07338_/X _13064_/Q _07339_/X vssd1 vssd1 vccd1 vccd1 _13064_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07277_ _11549_/X _07263_/X _13084_/Q _07264_/X vssd1 vssd1 vccd1 vccd1 _13084_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09016_ _09016_/A _09016_/B _11638_/X vssd1 vssd1 vccd1 vccd1 _12582_/D sky130_fd_sc_hd__and3_1
X_06228_ _06145_/X _06045_/A _06145_/X _06045_/A vssd1 vssd1 vccd1 vccd1 _06228_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_3_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06159_ _06025_/X _06158_/X _06025_/X _06158_/X vssd1 vssd1 vccd1 vccd1 _11963_/S
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_137_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09918_ _09914_/Y _09897_/X _06311_/A _09915_/X _09917_/X vssd1 vssd1 vccd1 vccd1
+ _09918_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09849_ _09849_/A vssd1 vssd1 vccd1 vccd1 _09849_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12860_ _12890_/CLK _12860_/D _08063_/X vssd1 vssd1 vccd1 vccd1 _12860_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11810_/X _12079_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12446_/D sky130_fd_sc_hd__mux2_1
XFILLER_2_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12872_/CLK _12791_/D _08389_/X vssd1 vssd1 vccd1 vccd1 _12791_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11741_/X _11369_/X _11774_/S vssd1 vssd1 vccd1 vccd1 _12425_/D sky130_fd_sc_hd__mux2_1
XPHY_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11387_/X _09184_/B _11675_/S vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10624_ _12415_/D _10610_/B _09428_/Y _12416_/D vssd1 vssd1 vccd1 vccd1 _10624_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10555_ _09333_/A _09333_/B _12362_/D vssd1 vssd1 vccd1 vccd1 _10555_/X sky130_fd_sc_hd__a21o_1
XFILLER_182_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ _13276_/CLK _13274_/D _06245_/X vssd1 vssd1 vccd1 vccd1 _13274_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10486_ _10486_/A vssd1 vssd1 vccd1 vccd1 _10486_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12225_ _06295_/Y _13158_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12156_ _10009_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12156_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11107_ _11107_/A vssd1 vssd1 vccd1 vccd1 _11107_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12087_ _10701_/Y _06634_/A _12758_/Q vssd1 vssd1 vccd1 vccd1 _12087_/X sky130_fd_sc_hd__mux2_2
XFILLER_110_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11038_ _12087_/X vssd1 vssd1 vccd1 vccd1 _11038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12989_ _12992_/CLK _12989_/D vssd1 vssd1 vccd1 vccd1 _12989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07200_ _07263_/A vssd1 vssd1 vccd1 vccd1 _07248_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08180_ _13128_/Q vssd1 vssd1 vccd1 vccd1 _08180_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07131_ _07161_/A vssd1 vssd1 vccd1 vccd1 _07131_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07062_ _07053_/X _07058_/X _06311_/Y _13155_/Q _07059_/X vssd1 vssd1 vccd1 vccd1
+ _13155_/D sky130_fd_sc_hd__a32o_1
XFILLER_118_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06013_ _09433_/A _09434_/B _11964_/S _09302_/A vssd1 vssd1 vccd1 vccd1 _09259_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_133_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07964_ _07985_/A vssd1 vssd1 vccd1 vccd1 _07964_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09703_ _06763_/Y _06768_/Y _09689_/Y _09690_/Y vssd1 vssd1 vccd1 vccd1 _09708_/A
+ sky130_fd_sc_hd__o22a_4
X_06915_ _06829_/X _06909_/Y _06769_/X _06914_/X vssd1 vssd1 vccd1 vccd1 _13185_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_96_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07895_ _07903_/A vssd1 vssd1 vccd1 vccd1 _07895_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09634_ _06865_/Y _06870_/Y _09617_/Y _09618_/Y vssd1 vssd1 vccd1 vccd1 _09640_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06846_ _12015_/X _06846_/B vssd1 vssd1 vccd1 vccd1 _06846_/X sky130_fd_sc_hd__or2_2
XFILLER_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09565_ _09572_/B vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__inv_2
X_06777_ _06806_/A vssd1 vssd1 vccd1 vccd1 _06777_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08516_ _08518_/A vssd1 vssd1 vccd1 vccd1 _08516_/X sky130_fd_sc_hd__clkbuf_1
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09496_ _09504_/A _09493_/Y _09495_/X vssd1 vssd1 vccd1 vccd1 _09496_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_130_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08447_ _13049_/Q vssd1 vssd1 vccd1 vccd1 _08447_/Y sky130_fd_sc_hd__inv_2
XPHY_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08378_ _12796_/Q _08374_/X _07287_/X _08375_/X vssd1 vssd1 vccd1 vccd1 _12796_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07329_ _11447_/X _07321_/X _13071_/Q _07324_/X vssd1 vssd1 vccd1 vccd1 _13071_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10340_ _12902_/Q vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__inv_2
XFILLER_87_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10271_ _09626_/Y _10166_/A _10270_/Y _10168_/A vssd1 vssd1 vccd1 vccd1 _10271_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12010_ _11090_/X _11081_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12010_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12912_ _12166_/X _12912_/D _07920_/X vssd1 vssd1 vccd1 vccd1 _12912_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12843_ _13146_/CLK _12843_/D _08249_/X vssd1 vssd1 vccd1 vccd1 _12843_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12774_ _12987_/CLK _12774_/D _08433_/X vssd1 vssd1 vccd1 vccd1 _12774_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _11724_/X _11915_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12441_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_48_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12458_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _10551_/Y _10550_/Y _11704_/S vssd1 vssd1 vccd1 vccd1 _12368_/D sky130_fd_sc_hd__mux2_1
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10607_ _10607_/A _11397_/X vssd1 vssd1 vccd1 vccd1 _10607_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_7_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11587_ _10426_/X _09183_/A _11592_/S vssd1 vssd1 vccd1 vccd1 _11587_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10538_ _09328_/A _09328_/B _09329_/B vssd1 vssd1 vccd1 vccd1 _10538_/X sky130_fd_sc_hd__a21bo_1
XFILLER_171_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13257_ _13257_/CLK _13257_/D _06338_/X vssd1 vssd1 vccd1 vccd1 _13257_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10469_ _10467_/B _10467_/C _10467_/A vssd1 vssd1 vccd1 vccd1 _10470_/C sky130_fd_sc_hd__o21a_1
XFILLER_97_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12208_ _12207_/X _12624_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12208_/X sky130_fd_sc_hd__mux2_1
X_13188_ _13190_/CLK _13188_/D _06885_/X vssd1 vssd1 vccd1 vccd1 _13188_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12139_ _12438_/Q _12138_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _12139_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06700_ _11986_/X _06698_/B _06698_/X vssd1 vssd1 vccd1 vccd1 _06700_/X sky130_fd_sc_hd__a21bo_1
X_07680_ _07680_/A vssd1 vssd1 vccd1 vccd1 _07726_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_64_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06631_ _11895_/X _06613_/X _11895_/X _06613_/X vssd1 vssd1 vccd1 vccd1 _06632_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09350_ _12408_/Q vssd1 vssd1 vccd1 vccd1 _09350_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06562_ _12174_/X _12173_/X vssd1 vssd1 vccd1 vccd1 _06562_/X sky130_fd_sc_hd__or2_1
X_08301_ _12827_/Q _11602_/X _08307_/S vssd1 vssd1 vccd1 vccd1 _12827_/D sky130_fd_sc_hd__mux2_1
XFILLER_166_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09281_ _08877_/X _07737_/X _07732_/X _12552_/Q _08908_/X vssd1 vssd1 vccd1 vccd1
+ _12552_/D sky130_fd_sc_hd__a41o_1
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06493_ _06427_/X _11077_/A _06356_/X _11086_/A _12195_/X vssd1 vssd1 vccd1 vccd1
+ _06494_/A sky130_fd_sc_hd__a221o_2
XFILLER_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08232_ _08232_/A _08232_/B _08232_/C _08231_/X vssd1 vssd1 vccd1 vccd1 _08238_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_21_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08163_ _08163_/A _08163_/B _08163_/C _08162_/X vssd1 vssd1 vccd1 vccd1 _08163_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_174_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07114_ _07176_/A vssd1 vssd1 vccd1 vccd1 _07177_/A sky130_fd_sc_hd__inv_2
XFILLER_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08094_ _08098_/A vssd1 vssd1 vccd1 vccd1 _08094_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07045_ _07037_/X _07040_/X _06278_/Y _13161_/Q _07042_/X vssd1 vssd1 vccd1 vccd1
+ _13161_/D sky130_fd_sc_hd__a32o_1
XFILLER_106_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08996_ _12593_/Q _11029_/A _12595_/Q _08996_/D vssd1 vssd1 vccd1 vccd1 _12597_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_125_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07947_ _07947_/A vssd1 vssd1 vccd1 vccd1 _08657_/A sky130_fd_sc_hd__buf_6
XFILLER_69_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07878_ _07803_/Y _07804_/X _13040_/Q _07809_/Y _07877_/Y vssd1 vssd1 vccd1 vccd1
+ _07879_/D sky130_fd_sc_hd__o221a_1
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09617_ _13191_/Q vssd1 vssd1 vccd1 vccd1 _09617_/Y sky130_fd_sc_hd__inv_2
X_06829_ _06887_/A vssd1 vssd1 vccd1 vccd1 _06829_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_141_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09548_ _09891_/A vssd1 vssd1 vccd1 vccd1 _09949_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ _13147_/Q _09475_/X _09476_/Y _09478_/X vssd1 vssd1 vccd1 vccd1 _09479_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11510_ _10394_/X _10794_/B _11513_/S vssd1 vssd1 vccd1 vccd1 _11510_/X sky130_fd_sc_hd__mux2_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12490_ _12490_/CLK _12490_/D vssd1 vssd1 vccd1 vccd1 _12490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11441_ _12916_/Q _09179_/C _11443_/S vssd1 vssd1 vccd1 vccd1 _11441_/X sky130_fd_sc_hd__mux2_1
XPHY_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11372_ _11371_/X _12426_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _11372_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13111_ _12167_/X _13111_/D _07209_/X vssd1 vssd1 vccd1 vccd1 _13111_/Q sky130_fd_sc_hd__dfrtp_1
X_10323_ _12894_/Q _12893_/Q _12895_/Q vssd1 vssd1 vccd1 vccd1 _10326_/B sky130_fd_sc_hd__and3_1
XFILLER_166_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13042_ _12165_/X _13042_/D _07400_/X vssd1 vssd1 vccd1 vccd1 _13042_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_124_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10254_ _13158_/Q vssd1 vssd1 vccd1 vccd1 _10254_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10185_ _12645_/Q vssd1 vssd1 vccd1 vccd1 _10185_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12826_ _12169_/X _12826_/D _08302_/X vssd1 vssd1 vccd1 vccd1 _12826_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12757_ _12769_/CLK _12757_/D _08528_/X vssd1 vssd1 vccd1 vccd1 _12757_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11707_/X _10629_/Y _11774_/S vssd1 vssd1 vccd1 vccd1 _12418_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12688_ _12688_/CLK _12688_/D _08732_/X vssd1 vssd1 vccd1 vccd1 _12688_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11639_ _10509_/X _12992_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11639_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08850_ _08849_/X _06300_/Y _08837_/X _12648_/Q vssd1 vssd1 vccd1 vccd1 _12648_/D
+ sky130_fd_sc_hd__o22a_1
X_07801_ _13035_/Q vssd1 vssd1 vccd1 vccd1 _07801_/Y sky130_fd_sc_hd__inv_2
X_08781_ _08781_/A vssd1 vssd1 vccd1 vccd1 _08781_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07732_ _09897_/A vssd1 vssd1 vccd1 vccd1 _07732_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07663_ _07663_/A vssd1 vssd1 vccd1 vccd1 _07668_/C sky130_fd_sc_hd__inv_2
XFILLER_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09402_ _09402_/A _09402_/B _09402_/C _09402_/D vssd1 vssd1 vccd1 vccd1 _09402_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06614_ _06611_/X _06612_/X _11895_/X _06613_/X vssd1 vssd1 vccd1 vccd1 _06614_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_197_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07594_ _12977_/Q vssd1 vssd1 vccd1 vccd1 _08977_/B sky130_fd_sc_hd__inv_2
XFILLER_53_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09333_ _09333_/A _09333_/B vssd1 vssd1 vccd1 vccd1 _12362_/D sky130_fd_sc_hd__nor2_1
X_06545_ _12176_/X _12175_/X _06539_/X _06540_/X _06544_/X vssd1 vssd1 vccd1 vccd1
+ _06546_/A sky130_fd_sc_hd__o32a_1
XFILLER_80_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09264_ _12941_/Q _09984_/A _09986_/B vssd1 vssd1 vccd1 vccd1 _09264_/X sky130_fd_sc_hd__and3_1
X_06476_ _09009_/A vssd1 vssd1 vccd1 vccd1 _06766_/A sky130_fd_sc_hd__buf_4
XFILLER_193_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ _13088_/Q _10420_/A _13096_/Q _10444_/B vssd1 vssd1 vccd1 vccd1 _08215_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09195_ _12490_/Q _09190_/X _09180_/A _09192_/X vssd1 vssd1 vccd1 vccd1 _12490_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08146_ _12823_/Q vssd1 vssd1 vccd1 vccd1 _10454_/A sky130_fd_sc_hd__inv_2
XFILLER_174_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08077_ _08085_/A vssd1 vssd1 vccd1 vccd1 _08077_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07028_ _06663_/X _12181_/X _06415_/B _13165_/Q vssd1 vssd1 vccd1 vccd1 _13165_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput304 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _07101_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput315 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _07096_/C sky130_fd_sc_hd__clkbuf_1
Xinput326 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 input326/X sky130_fd_sc_hd__buf_1
XFILLER_103_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput337 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 input337/X sky130_fd_sc_hd__buf_2
X_08979_ _13006_/Q _13005_/Q _11147_/A vssd1 vssd1 vccd1 vccd1 _12603_/D sky130_fd_sc_hd__o21a_1
Xinput348 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 _10794_/C sky130_fd_sc_hd__buf_6
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput359 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 _09183_/A sky130_fd_sc_hd__buf_8
XFILLER_75_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11990_ _11123_/X _11116_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _11990_/X sky130_fd_sc_hd__mux2_2
XFILLER_21_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10941_ _12533_/Q _12345_/Q _12533_/Q _12345_/Q vssd1 vssd1 vccd1 vccd1 _10945_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10872_ _12335_/Q vssd1 vssd1 vccd1 vccd1 _10873_/B sky130_fd_sc_hd__inv_2
XFILLER_72_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _12688_/CLK _12612_/Q _08967_/X vssd1 vssd1 vccd1 vccd1 _12611_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12542_ _12547_/CLK _12542_/D vssd1 vssd1 vccd1 vccd1 _12542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12473_ _12474_/CLK _12473_/D vssd1 vssd1 vccd1 vccd1 _12473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11424_ _12899_/Q _09184_/B _11433_/S vssd1 vssd1 vccd1 vccd1 _11424_/X sky130_fd_sc_hd__mux2_1
X_11355_ _09465_/X _12992_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _12319_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10306_ _09934_/Y _09968_/X _10297_/X _10305_/X vssd1 vssd1 vccd1 vccd1 _10306_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_140_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11286_ vssd1 vssd1 vccd1 vccd1 _11286_/HI _11286_/LO sky130_fd_sc_hd__conb_1
XFILLER_134_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13025_ _12164_/X _13025_/D _07452_/X vssd1 vssd1 vccd1 vccd1 _13025_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_156_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10237_ _12887_/Q vssd1 vssd1 vccd1 vccd1 _10237_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10168_ _10168_/A vssd1 vssd1 vccd1 vccd1 _10168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_187_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10099_ _12641_/Q vssd1 vssd1 vccd1 vccd1 _10099_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_wb_clk_i _12960_/CLK vssd1 vssd1 vccd1 vccd1 _12509_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12809_ _12169_/X _12809_/D _08342_/X vssd1 vssd1 vccd1 vccd1 _12809_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06330_ _06112_/Y _06113_/Y _06125_/C _06125_/B vssd1 vssd1 vccd1 vccd1 _06330_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06261_ _06258_/Y _06247_/X _06217_/A _06260_/X vssd1 vssd1 vccd1 vccd1 _13272_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_198_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08000_ _08004_/A vssd1 vssd1 vccd1 vccd1 _08000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06192_ _06035_/B _06186_/X _06035_/B _06186_/X vssd1 vssd1 vccd1 vccd1 _06192_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_156_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09951_ _08777_/Y _09943_/X _06237_/X _09949_/X _09950_/X vssd1 vssd1 vccd1 vccd1
+ _09951_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_132_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08902_ _08898_/X _06323_/Y _08893_/X _12628_/Q vssd1 vssd1 vccd1 vccd1 _12628_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_98_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09882_ _09873_/Y _09874_/X _09857_/Y _09880_/B vssd1 vssd1 vccd1 vccd1 _09882_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_83_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08833_ _08814_/A _08781_/A _06346_/Y _12655_/Q _08567_/A vssd1 vssd1 vccd1 vccd1
+ _12655_/D sky130_fd_sc_hd__a32o_1
XFILLER_44_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08764_ _08764_/A vssd1 vssd1 vccd1 vccd1 _08764_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ _12953_/Q _07707_/X _12952_/Q _07705_/X _07714_/X vssd1 vssd1 vccd1 vccd1
+ _12953_/D sky130_fd_sc_hd__o221a_1
XFILLER_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08695_ _08699_/A vssd1 vssd1 vccd1 vccd1 _08695_/X sky130_fd_sc_hd__clkbuf_1
XPHY_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07646_ _12961_/Q _12960_/Q _07660_/C _07646_/D vssd1 vssd1 vccd1 vccd1 _07652_/A
+ sky130_fd_sc_hd__or4_4
XPHY_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07577_ _12985_/Q _07574_/X _09185_/A _07575_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _12985_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ _09316_/A vssd1 vssd1 vccd1 vccd1 _12091_/S sky130_fd_sc_hd__clkinv_4
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06528_ _12621_/Q vssd1 vssd1 vccd1 vccd1 _06528_/X sky130_fd_sc_hd__buf_2
XFILLER_90_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09247_ _09247_/A _11691_/S vssd1 vssd1 vccd1 vccd1 _09250_/A sky130_fd_sc_hd__nand2_1
XFILLER_142_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06459_ _06769_/A vssd1 vssd1 vccd1 vccd1 _06459_/X sky130_fd_sc_hd__buf_2
XFILLER_5_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09178_ _12468_/Q _09304_/B vssd1 vssd1 vccd1 vccd1 _10655_/B sky130_fd_sc_hd__or2_4
XFILLER_135_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ _13123_/Q vssd1 vssd1 vccd1 vccd1 _08129_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11140_ _10773_/A _10737_/A _13246_/Q _10738_/X _10739_/X vssd1 vssd1 vccd1 vccd1
+ _11140_/X sky130_fd_sc_hd__a221o_1
XFILLER_122_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11071_ _11071_/A vssd1 vssd1 vccd1 vccd1 _11071_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput101 la_data_in[40] vssd1 vssd1 vccd1 vccd1 input101/X sky130_fd_sc_hd__buf_1
XFILLER_131_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput112 la_data_in[50] vssd1 vssd1 vccd1 vccd1 input112/X sky130_fd_sc_hd__buf_1
X_10022_ _13147_/Q vssd1 vssd1 vccd1 vccd1 _10022_/Y sky130_fd_sc_hd__inv_2
Xinput123 la_data_in[60] vssd1 vssd1 vccd1 vccd1 input123/X sky130_fd_sc_hd__buf_1
Xinput134 la_data_in[70] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__buf_1
XFILLER_130_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput145 la_data_in[80] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_hd__buf_1
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput156 la_data_in[90] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__buf_1
Xinput167 la_oenb[0] vssd1 vssd1 vccd1 vccd1 _11344_/A sky130_fd_sc_hd__buf_4
Xinput178 la_oenb[10] vssd1 vssd1 vccd1 vccd1 input178/X sky130_fd_sc_hd__buf_1
XFILLER_64_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput189 la_oenb[11] vssd1 vssd1 vccd1 vccd1 input189/X sky130_fd_sc_hd__buf_1
XFILLER_45_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11973_ _10068_/Y _12789_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11973_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10924_ _12527_/Q _12339_/Q _10923_/X _10908_/X _10915_/A vssd1 vssd1 vccd1 vccd1
+ _10924_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_17_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10855_ _12333_/Q vssd1 vssd1 vccd1 vccd1 _10855_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _10755_/X _10731_/X _06371_/X _10732_/X _10733_/X vssd1 vssd1 vccd1 vccd1
+ _10786_/X sky130_fd_sc_hd__a221o_1
XFILLER_197_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12525_ _12535_/CLK _12525_/D vssd1 vssd1 vccd1 vccd1 _12525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12456_ _12458_/CLK _12456_/D vssd1 vssd1 vccd1 vccd1 _12456_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_110_wb_clk_i clkbuf_opt_3_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12743_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11407_ _11040_/X _10746_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _11407_/X sky130_fd_sc_hd__mux2_1
X_12387_ _12492_/CLK _12387_/D vssd1 vssd1 vccd1 vccd1 _12409_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11338_ vssd1 vssd1 vccd1 vccd1 _11338_/HI _11338_/LO sky130_fd_sc_hd__conb_1
XFILLER_180_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11269_ vssd1 vssd1 vccd1 vccd1 _11269_/HI _11269_/LO sky130_fd_sc_hd__conb_1
XFILLER_122_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13008_ _13008_/CLK _13008_/D vssd1 vssd1 vccd1 vccd1 _13008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07500_ _13008_/Q vssd1 vssd1 vccd1 vccd1 _09279_/C sky130_fd_sc_hd__inv_2
X_08480_ _13058_/Q _10362_/B vssd1 vssd1 vccd1 vccd1 _08480_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07431_ _11475_/X _07429_/X _13034_/Q _07430_/X vssd1 vssd1 vccd1 vccd1 _13034_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07362_ _07362_/A vssd1 vssd1 vccd1 vccd1 _07375_/A sky130_fd_sc_hd__buf_2
XFILLER_50_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09101_ _12535_/Q _09099_/X _10792_/A _09100_/X vssd1 vssd1 vccd1 vccd1 _12535_/D
+ sky130_fd_sc_hd__a22o_1
X_06313_ _06313_/A vssd1 vssd1 vccd1 vccd1 _06313_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07293_ _09185_/B vssd1 vssd1 vccd1 vccd1 _07293_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_149_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09032_ _12180_/X _09288_/A vssd1 vssd1 vccd1 vccd1 _12573_/D sky130_fd_sc_hd__and2_1
XFILLER_136_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06244_ _06240_/Y _06216_/X _06217_/X _06243_/X vssd1 vssd1 vccd1 vccd1 _13275_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_50_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06175_ _06175_/A _06175_/B vssd1 vssd1 vccd1 vccd1 _06320_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09934_ _12668_/Q vssd1 vssd1 vccd1 vccd1 _09934_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09865_ _13238_/Q _09864_/A _09686_/X _09864_/Y vssd1 vssd1 vccd1 vccd1 _09879_/A
+ sky130_fd_sc_hd__a22o_1
X_08816_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08816_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09796_ _09886_/A _09796_/B vssd1 vssd1 vccd1 vccd1 _09796_/X sky130_fd_sc_hd__or2_1
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08747_ _08747_/A vssd1 vssd1 vccd1 vccd1 _08747_/X sky130_fd_sc_hd__clkbuf_1
XPHY_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08678_/X sky130_fd_sc_hd__clkbuf_1
XPHY_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07629_ _07661_/A _12953_/Q _07658_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07670_/C
+ sky130_fd_sc_hd__or4_4
XPHY_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _12421_/Q _10636_/Y _08929_/B vssd1 vssd1 vccd1 vccd1 _10640_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10571_ _12399_/D _10570_/A _12400_/D vssd1 vssd1 vccd1 vccd1 _10571_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_167_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12310_ _12951_/CLK _12310_/D vssd1 vssd1 vccd1 vccd1 _12310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12241_ _12775_/Q _12848_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12241_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12172_ _11141_/X _11136_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12172_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11123_ _10742_/X _11054_/A _13251_/Q _11055_/A _11899_/X vssd1 vssd1 vccd1 vccd1
+ _11123_/X sky130_fd_sc_hd__a221o_1
XFILLER_174_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11054_ _11054_/A vssd1 vssd1 vccd1 vccd1 _11054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10005_ _08767_/Y _10003_/X _06222_/Y _10000_/X _10001_/X vssd1 vssd1 vccd1 vccd1
+ _10005_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11956_ _09872_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11956_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ _12340_/Q vssd1 vssd1 vccd1 vccd1 _10907_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11887_ _10623_/X _12415_/D _11889_/S vssd1 vssd1 vccd1 vccd1 _11887_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10838_ _12330_/Q vssd1 vssd1 vccd1 vccd1 _10838_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10769_ _11107_/A vssd1 vssd1 vccd1 vccd1 _10769_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12508_ _12509_/CLK _12508_/D vssd1 vssd1 vccd1 vccd1 _12508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12439_ _12485_/CLK _12439_/D vssd1 vssd1 vccd1 vccd1 _12439_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput405 _11182_/LO vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput416 _11183_/LO vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput427 _11184_/LO vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput438 _11347_/X vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput449 _11318_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07980_ _07980_/A vssd1 vssd1 vccd1 vccd1 _07980_/X sky130_fd_sc_hd__buf_2
XFILLER_113_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06931_ _06931_/A vssd1 vssd1 vccd1 vccd1 _06935_/A sky130_fd_sc_hd__inv_2
XFILLER_45_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09650_ _09635_/Y _06844_/Y _09637_/Y _09638_/Y vssd1 vssd1 vccd1 vccd1 _09655_/A
+ sky130_fd_sc_hd__o22a_1
X_06862_ _06719_/X _06810_/Y _06861_/X _06841_/X _13191_/Q vssd1 vssd1 vccd1 vccd1
+ _13191_/D sky130_fd_sc_hd__a32o_1
X_08601_ _11949_/X _08592_/X _12740_/Q _08593_/X vssd1 vssd1 vccd1 vccd1 _12740_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09581_ _09607_/A vssd1 vssd1 vccd1 vccd1 _09582_/B sky130_fd_sc_hd__inv_2
XFILLER_83_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06793_ _06658_/A _06783_/X _06791_/X _06646_/X _06792_/Y vssd1 vssd1 vccd1 vccd1
+ _06794_/A sky130_fd_sc_hd__a32o_1
XFILLER_94_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08532_ _08519_/X _12238_/X _06396_/A _10701_/A vssd1 vssd1 vccd1 vccd1 _12756_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08463_ _13057_/Q _10357_/A _13070_/Q _10393_/A vssd1 vssd1 vccd1 vccd1 _08467_/B
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07414_ _07475_/A vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_196_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08394_ _12789_/Q _08374_/A _07309_/X _08375_/A vssd1 vssd1 vccd1 vccd1 _12789_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07345_ _07345_/A vssd1 vssd1 vccd1 vccd1 _07345_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07276_ _07280_/A vssd1 vssd1 vccd1 vccd1 _07276_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09015_ _09016_/A _09016_/B _11639_/X vssd1 vssd1 vccd1 vccd1 _12583_/D sky130_fd_sc_hd__and3_1
X_06227_ _13278_/Q vssd1 vssd1 vccd1 vccd1 _06227_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06158_ _06185_/A _06035_/X _06197_/B _06145_/X _06157_/Y vssd1 vssd1 vccd1 vccd1
+ _06158_/X sky130_fd_sc_hd__o41a_1
XFILLER_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06089_ _06087_/Y _06088_/Y _12727_/Q _12695_/Q vssd1 vssd1 vccd1 vccd1 _06090_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09917_ _12885_/Q _09935_/B vssd1 vssd1 vccd1 vccd1 _09917_/X sky130_fd_sc_hd__or2_1
XFILLER_144_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09848_ _09848_/A _09868_/A vssd1 vssd1 vccd1 vccd1 _09851_/B sky130_fd_sc_hd__or2_1
XFILLER_46_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09779_/A _09779_/B vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__or2_1
XPHY_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _12079_/X _11809_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11810_/X sky130_fd_sc_hd__mux2_1
XPHY_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12840_/CLK _12790_/D _08391_/X vssd1 vssd1 vccd1 vccd1 _12790_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_199_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11741_ _11369_/X _11740_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11741_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11671_/X _11389_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12378_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _12415_/D _10615_/B _09428_/Y _11888_/S _11406_/X vssd1 vssd1 vccd1 vccd1
+ _10623_/X sky130_fd_sc_hd__o221a_1
XFILLER_23_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ _11393_/X _10554_/B vssd1 vssd1 vccd1 vccd1 _10554_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13273_ _13276_/CLK _13273_/D _06251_/X vssd1 vssd1 vccd1 vccd1 _13273_/Q sky130_fd_sc_hd__dfrtp_1
X_10485_ _10484_/A _10484_/B _10459_/X _10486_/A vssd1 vssd1 vccd1 vccd1 _10485_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12224_ _12223_/X _12632_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12224_/X sky130_fd_sc_hd__mux2_2
XFILLER_135_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12155_ _10008_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12155_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11106_ _10779_/X _11077_/X _13245_/Q _11086_/X _11087_/X vssd1 vssd1 vccd1 vccd1
+ _11106_/X sky130_fd_sc_hd__a221o_1
XFILLER_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12086_ _12085_/X _12447_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12086_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11037_ _11071_/A vssd1 vssd1 vccd1 vccd1 _11037_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12988_ _12992_/CLK _12988_/D vssd1 vssd1 vccd1 vccd1 _12988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11939_ _09628_/X _12800_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11939_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07130_ _07160_/A vssd1 vssd1 vccd1 vccd1 _07130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07061_ _07063_/A vssd1 vssd1 vccd1 vccd1 _07061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06012_ _11966_/S vssd1 vssd1 vccd1 vccd1 _09302_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07963_ _08038_/A vssd1 vssd1 vccd1 vccd1 _07985_/A sky130_fd_sc_hd__buf_2
XFILLER_141_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09702_ _09687_/X _09691_/X _09686_/X _09692_/X vssd1 vssd1 vccd1 vccd1 _09711_/A
+ sky130_fd_sc_hd__o22a_2
X_06914_ _06910_/X _06911_/X _06904_/X _06896_/X _06913_/X vssd1 vssd1 vccd1 vccd1
+ _06914_/X sky130_fd_sc_hd__o221a_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07894_ _12924_/Q _11513_/X _07904_/S vssd1 vssd1 vccd1 vccd1 _12924_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06845_ _12011_/X vssd1 vssd1 vccd1 vccd1 _06846_/B sky130_fd_sc_hd__inv_2
XFILLER_28_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09633_ _09608_/Y _09632_/B _09675_/A _09632_/X vssd1 vssd1 vccd1 vccd1 _09714_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09564_ _09550_/A _09550_/B _09563_/A _09550_/Y _09563_/Y vssd1 vssd1 vccd1 vccd1
+ _09572_/B sky130_fd_sc_hd__o32a_1
X_06776_ _06658_/X _06768_/Y _06769_/X _06775_/X vssd1 vssd1 vccd1 vccd1 _13201_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08515_ _08504_/X _12252_/X _08514_/X _12763_/Q vssd1 vssd1 vccd1 vccd1 _12763_/D
+ sky130_fd_sc_hd__o22a_1
X_09495_ _13149_/Q _07737_/A _09494_/Y _09478_/X vssd1 vssd1 vccd1 vccd1 _09495_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08446_ _13068_/Q vssd1 vssd1 vccd1 vccd1 _08446_/Y sky130_fd_sc_hd__inv_2
XPHY_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08377_ _08385_/A vssd1 vssd1 vccd1 vccd1 _08377_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_196_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07328_ _07330_/A vssd1 vssd1 vccd1 vccd1 _07328_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07259_ _11556_/X _07248_/X _13091_/Q _07249_/X vssd1 vssd1 vccd1 vccd1 _13091_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10270_ _12650_/Q vssd1 vssd1 vccd1 vccd1 _10270_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12911_ _12166_/X _12911_/D _07923_/X vssd1 vssd1 vccd1 vccd1 _12911_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_150_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12842_ _13146_/CLK _12842_/D _08253_/X vssd1 vssd1 vccd1 vccd1 _12842_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12773_/CLK _12773_/D _08436_/X vssd1 vssd1 vccd1 vccd1 _12773_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11724_ _11915_/X _11723_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11724_/X sky130_fd_sc_hd__mux2_1
XPHY_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11655_ _10547_/Y _10546_/Y _11704_/S vssd1 vssd1 vccd1 vccd1 _12367_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10606_ _12409_/D _09385_/Y _10602_/Y _12410_/D _10603_/X vssd1 vssd1 vccd1 vccd1
+ _10606_/X sky130_fd_sc_hd__a32o_1
XPHY_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_88_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _12646_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11586_ _10423_/X _09185_/A _11592_/S vssd1 vssd1 vccd1 vccd1 _11586_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10537_ _11361_/X _10554_/B vssd1 vssd1 vccd1 vccd1 _10537_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_17_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12485_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13256_ _13256_/CLK _13256_/D _06344_/X vssd1 vssd1 vccd1 vccd1 _13256_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ _10468_/A vssd1 vssd1 vccd1 vccd1 _10472_/C sky130_fd_sc_hd__inv_2
XFILLER_124_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12207_ _06342_/Y _13149_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12207_/X sky130_fd_sc_hd__mux2_1
X_13187_ _13190_/CLK _13187_/D _06889_/X vssd1 vssd1 vccd1 vccd1 _13187_/Q sky130_fd_sc_hd__dfrtp_1
X_10399_ _10399_/A vssd1 vssd1 vccd1 vccd1 _10399_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12138_ _10676_/X _08952_/B _12138_/S vssd1 vssd1 vccd1 vccd1 _12138_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12069_ _12445_/Q _12068_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06630_ _12621_/Q vssd1 vssd1 vccd1 vccd1 _06630_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06561_ _13222_/Q vssd1 vssd1 vccd1 vccd1 _09798_/B sky130_fd_sc_hd__inv_2
X_08300_ _08311_/A vssd1 vssd1 vccd1 vccd1 _08300_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09280_ _07726_/A _09278_/Y _09279_/X vssd1 vssd1 vccd1 vccd1 _12311_/D sky130_fd_sc_hd__o21ai_1
X_06492_ _11077_/A vssd1 vssd1 vccd1 vccd1 _11086_/A sky130_fd_sc_hd__inv_2
XFILLER_20_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08231_ _13096_/Q _10444_/B _13110_/Q _10480_/A vssd1 vssd1 vccd1 vccd1 _08231_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08162_ _08153_/X _08162_/B _08162_/C _08162_/D vssd1 vssd1 vccd1 vccd1 _08162_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_158_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07113_ _07160_/A vssd1 vssd1 vccd1 vccd1 _07113_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08093_ _12850_/Q _08082_/X _07293_/X _08083_/X vssd1 vssd1 vccd1 vccd1 _12850_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07044_ _07046_/A vssd1 vssd1 vccd1 vccd1 _07044_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_173_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08995_ _08996_/D _11029_/A _08995_/C _12593_/Q vssd1 vssd1 vccd1 vccd1 _12598_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07946_ _07821_/X _11490_/X _07946_/S vssd1 vssd1 vccd1 vccd1 _12901_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07877_ _13025_/Q _10368_/B vssd1 vssd1 vccd1 vccd1 _07877_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09616_ _13190_/Q _13189_/Q _06865_/Y _06870_/Y vssd1 vssd1 vccd1 vccd1 _09618_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06828_ _06863_/A vssd1 vssd1 vccd1 vccd1 _06828_/X sky130_fd_sc_hd__buf_1
XFILLER_3_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06759_ _12002_/X _11999_/X _12002_/X _11999_/X vssd1 vssd1 vccd1 vccd1 _06759_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09547_ _09547_/A vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__inv_2
XFILLER_110_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ _09939_/B vssd1 vssd1 vccd1 vccd1 _09478_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12726_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_08429_ _08433_/A vssd1 vssd1 vccd1 vccd1 _08429_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11440_ _12915_/Q _09179_/D _11443_/S vssd1 vssd1 vccd1 vccd1 _11440_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11371_ _11370_/X _12426_/Q _12103_/S vssd1 vssd1 vccd1 vccd1 _11371_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10322_ _10318_/Y _07822_/Y _07823_/Y vssd1 vssd1 vccd1 vccd1 _10325_/A sky130_fd_sc_hd__o21a_1
XFILLER_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13110_ _12167_/X _13110_/D _07211_/X vssd1 vssd1 vccd1 vccd1 _13110_/Q sky130_fd_sc_hd__dfrtp_1
X_13041_ _12166_/A0 _13041_/D _07402_/X vssd1 vssd1 vccd1 vccd1 _13146_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_106_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10253_ _12633_/Q vssd1 vssd1 vccd1 vccd1 _10253_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10184_ _13154_/Q vssd1 vssd1 vccd1 vccd1 _10184_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_135_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13159_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12825_ _12169_/X _12825_/D _08304_/X vssd1 vssd1 vccd1 vccd1 _12825_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _13241_/CLK _12756_/D _08530_/X vssd1 vssd1 vccd1 vccd1 _12756_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11707_ _10629_/Y _10632_/Y _11818_/S vssd1 vssd1 vccd1 vccd1 _11707_/X sky130_fd_sc_hd__mux2_1
XPHY_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _12719_/CLK _12687_/D _08734_/X vssd1 vssd1 vccd1 vccd1 _12687_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11638_ _10508_/X _12991_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11638_/X sky130_fd_sc_hd__mux2_1
XPHY_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11569_ _12826_/Q _09179_/D _11569_/S vssd1 vssd1 vccd1 vccd1 _11569_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13239_ _13241_/CLK _13239_/D _06409_/X vssd1 vssd1 vccd1 vccd1 _13239_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_171_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07800_ _12896_/Q vssd1 vssd1 vccd1 vccd1 _07800_/X sky130_fd_sc_hd__clkbuf_2
X_08780_ _12674_/Q vssd1 vssd1 vccd1 vccd1 _08780_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07731_ _09546_/A vssd1 vssd1 vccd1 vccd1 _09897_/A sky130_fd_sc_hd__buf_2
XFILLER_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07662_ _12960_/Q _07688_/A _07661_/C _07689_/C _07652_/X vssd1 vssd1 vccd1 vccd1
+ _07663_/A sky130_fd_sc_hd__o311a_1
XFILLER_53_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09401_ _12462_/Q _10562_/A _12545_/Q _09399_/Y _09400_/X vssd1 vssd1 vccd1 vccd1
+ _09402_/D sky130_fd_sc_hd__o221a_1
X_06613_ _06611_/X _06612_/X _06611_/X _06612_/X vssd1 vssd1 vccd1 vccd1 _06613_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07593_ _09268_/B vssd1 vssd1 vccd1 vccd1 _09288_/A sky130_fd_sc_hd__buf_2
XFILLER_129_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09332_ _09332_/A _10548_/A vssd1 vssd1 vccd1 vccd1 _09333_/B sky130_fd_sc_hd__or2_1
XFILLER_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06544_ _06541_/X _06542_/X _12179_/X _06543_/X vssd1 vssd1 vccd1 vccd1 _06544_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09263_ _10015_/B _09029_/B _09283_/A _09262_/X vssd1 vssd1 vccd1 vccd1 _12303_/D
+ sky130_fd_sc_hd__o31ai_1
X_06475_ _06440_/X _06466_/Y _06420_/X _06474_/X vssd1 vssd1 vccd1 vccd1 _13232_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_166_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08214_ _12821_/Q vssd1 vssd1 vccd1 vccd1 _10455_/A sky130_fd_sc_hd__inv_2
XFILLER_14_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09194_ _12491_/Q _09190_/X _09179_/D _09192_/X vssd1 vssd1 vccd1 vccd1 _12491_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08145_ _13129_/Q _10444_/A _13142_/Q _10480_/A vssd1 vssd1 vccd1 vccd1 _08151_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08076_ _12857_/Q _08066_/X _07986_/X _08068_/X vssd1 vssd1 vccd1 vccd1 _12857_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07027_ _07046_/A vssd1 vssd1 vccd1 vccd1 _07027_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput305 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _07101_/D sky130_fd_sc_hd__clkbuf_1
Xinput316 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 _07100_/A sky130_fd_sc_hd__clkbuf_1
Xinput327 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 input327/X sky130_fd_sc_hd__buf_1
Xinput338 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 input338/X sky130_fd_sc_hd__buf_2
XFILLER_103_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput349 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 _10794_/B sky130_fd_sc_hd__buf_4
X_08978_ _08978_/A vssd1 vssd1 vccd1 vccd1 _11147_/A sky130_fd_sc_hd__buf_6
XFILLER_102_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07929_ _07931_/A vssd1 vssd1 vccd1 vccd1 _07929_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10940_ _10945_/C _10939_/Y _10945_/C _10939_/Y vssd1 vssd1 vccd1 vccd1 _12344_/D
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_1_wb_clk_i clkbuf_2_1_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10871_ _12523_/Q vssd1 vssd1 vccd1 vccd1 _10873_/A sky130_fd_sc_hd__inv_2
XFILLER_25_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _13268_/CLK _12611_/Q _08968_/X vssd1 vssd1 vccd1 vccd1 _12610_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _12541_/CLK _12541_/D vssd1 vssd1 vccd1 vccd1 _12541_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12472_ _12472_/CLK _12472_/D vssd1 vssd1 vccd1 vccd1 _12472_/Q sky130_fd_sc_hd__dfxtp_1
X_11423_ _12898_/Q input356/X _11433_/S vssd1 vssd1 vccd1 vccd1 _11423_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11354_ _09462_/X _12991_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _12318_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10305_ _10298_/Y _10038_/X _09649_/Y _10033_/X _10304_/X vssd1 vssd1 vccd1 vccd1
+ _10305_/X sky130_fd_sc_hd__o221a_1
X_11285_ vssd1 vssd1 vccd1 vccd1 _11285_/HI _11285_/LO sky130_fd_sc_hd__conb_1
XFILLER_113_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13024_ _12164_/X _13024_/D _07454_/X vssd1 vssd1 vccd1 vccd1 _13024_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10236_ _12871_/Q vssd1 vssd1 vccd1 vccd1 _10236_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10167_ _12644_/Q vssd1 vssd1 vccd1 vccd1 _10167_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10098_ _13150_/Q vssd1 vssd1 vccd1 vccd1 _10098_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ _12169_/X _12808_/D _08344_/X vssd1 vssd1 vccd1 vccd1 _12808_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_32_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12471_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12739_ _12743_/CLK _12739_/D _08602_/X vssd1 vssd1 vccd1 vccd1 _12739_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_187_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06260_ _06259_/A _06253_/Y _06259_/Y _06253_/A vssd1 vssd1 vccd1 vccd1 _06260_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_124_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06191_ _13284_/Q vssd1 vssd1 vccd1 vccd1 _06191_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09950_ _09950_/A vssd1 vssd1 vccd1 vccd1 _09950_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08901_ _08912_/A vssd1 vssd1 vccd1 vccd1 _08901_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09881_ _09881_/A _09881_/B vssd1 vssd1 vccd1 vccd1 _09881_/X sky130_fd_sc_hd__or2_1
XFILLER_97_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08832_ _08836_/A vssd1 vssd1 vccd1 vccd1 _08832_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08763_ _12679_/Q vssd1 vssd1 vccd1 vccd1 _08763_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07714_ _09268_/B vssd1 vssd1 vccd1 vccd1 _07714_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _11838_/X _08685_/X _12704_/Q _08686_/X vssd1 vssd1 vccd1 vccd1 _12704_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07645_ _07659_/A _07689_/B vssd1 vssd1 vccd1 vccd1 _07648_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07576_ _08978_/A vssd1 vssd1 vccd1 vccd1 _07576_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09315_ _09315_/A vssd1 vssd1 vccd1 vccd1 _12138_/S sky130_fd_sc_hd__inv_2
X_06527_ _06527_/A _06527_/B vssd1 vssd1 vccd1 vccd1 _06527_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09246_ _09246_/A vssd1 vssd1 vccd1 vccd1 _11691_/S sky130_fd_sc_hd__buf_4
XFILLER_22_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06458_ _06458_/A _06458_/B vssd1 vssd1 vccd1 vccd1 _06458_/X sky130_fd_sc_hd__or2_1
XFILLER_182_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09177_ _09437_/A _10527_/D vssd1 vssd1 vccd1 vccd1 _09304_/B sky130_fd_sc_hd__or2_2
XFILLER_119_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06389_ _13245_/Q vssd1 vssd1 vccd1 vccd1 _06389_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_175_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08128_ _12825_/Q vssd1 vssd1 vccd1 vccd1 _08128_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08059_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08059_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11070_ _06376_/X _11045_/X _08535_/A _10758_/X _07030_/X vssd1 vssd1 vccd1 vccd1
+ _11070_/X sky130_fd_sc_hd__a32o_1
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput102 la_data_in[41] vssd1 vssd1 vccd1 vccd1 input102/X sky130_fd_sc_hd__buf_1
X_10021_ _10017_/Y _10018_/X _10019_/Y _10020_/X vssd1 vssd1 vccd1 vccd1 _10041_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_103_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput113 la_data_in[51] vssd1 vssd1 vccd1 vccd1 input113/X sky130_fd_sc_hd__buf_1
XFILLER_62_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput124 la_data_in[61] vssd1 vssd1 vccd1 vccd1 input124/X sky130_fd_sc_hd__buf_1
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput135 la_data_in[71] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_hd__buf_1
XFILLER_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput146 la_data_in[81] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_hd__buf_1
Xinput157 la_data_in[91] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_hd__buf_1
Xinput168 la_oenb[100] vssd1 vssd1 vccd1 vccd1 input168/X sky130_fd_sc_hd__buf_1
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput179 la_oenb[110] vssd1 vssd1 vccd1 vccd1 input179/X sky130_fd_sc_hd__buf_1
XFILLER_56_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11972_ _10041_/Y _12788_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11972_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10923_ _12526_/Q _12338_/Q _10900_/Y vssd1 vssd1 vccd1 vccd1 _10923_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10854_ _12521_/Q vssd1 vssd1 vccd1 vccd1 _10854_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10785_ _10742_/X _10731_/X _06368_/X _10732_/X _10733_/X vssd1 vssd1 vccd1 vccd1
+ _10785_/X sky130_fd_sc_hd__a221o_1
XFILLER_200_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12524_ _12535_/CLK _12524_/D vssd1 vssd1 vccd1 vccd1 _12524_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12455_ _12455_/CLK _12455_/D vssd1 vssd1 vccd1 vccd1 _12455_/Q sky130_fd_sc_hd__dfxtp_1
X_11406_ _10619_/B _10610_/B _11406_/S vssd1 vssd1 vccd1 vccd1 _11406_/X sky130_fd_sc_hd__mux2_1
X_12386_ _12467_/CLK _12386_/D vssd1 vssd1 vccd1 vccd1 _12408_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_126_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11337_ vssd1 vssd1 vccd1 vccd1 _11337_/HI _11337_/LO sky130_fd_sc_hd__conb_1
XFILLER_67_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_150_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12890_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ vssd1 vssd1 vccd1 vccd1 _11268_/HI _11268_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _13008_/CLK _13007_/D vssd1 vssd1 vccd1 vccd1 _13007_/Q sky130_fd_sc_hd__dfxtp_1
X_10219_ _12886_/Q vssd1 vssd1 vccd1 vccd1 _10219_/Y sky130_fd_sc_hd__inv_2
X_11199_ vssd1 vssd1 vccd1 vccd1 _11199_/HI _11199_/LO sky130_fd_sc_hd__conb_1
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07430_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07430_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07361_ _11434_/X _07353_/X _13058_/Q _07354_/X vssd1 vssd1 vccd1 vccd1 _13058_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09100_ _09116_/A vssd1 vssd1 vccd1 vccd1 _09100_/X sky130_fd_sc_hd__clkbuf_2
X_06312_ _06303_/X _06281_/X _06311_/Y _13263_/Q _06306_/X vssd1 vssd1 vccd1 vccd1
+ _13263_/D sky130_fd_sc_hd__a32o_1
XFILLER_149_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07292_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07292_/X sky130_fd_sc_hd__clkbuf_1
X_09031_ _09027_/Y _09030_/Y _07695_/X vssd1 vssd1 vccd1 vccd1 _12574_/D sky130_fd_sc_hd__o21a_1
X_06243_ _06056_/A _06242_/Y _06056_/A _06242_/Y vssd1 vssd1 vccd1 vccd1 _06243_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_175_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06174_ _06174_/A vssd1 vssd1 vccd1 vccd1 _06174_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09933_ _09931_/Y _09922_/X _06283_/A _09915_/X _09932_/X vssd1 vssd1 vccd1 vccd1
+ _09933_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09864_ _09864_/A vssd1 vssd1 vccd1 vccd1 _09864_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08815_ _08814_/X _08801_/X _06305_/X _12663_/Q _08811_/X vssd1 vssd1 vccd1 vccd1
+ _12663_/D sky130_fd_sc_hd__a32o_1
XFILLER_100_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09795_ _09802_/B _09794_/Y _09792_/A _09794_/A _09492_/A vssd1 vssd1 vccd1 vccd1
+ _09796_/B sky130_fd_sc_hd__o221a_1
XFILLER_61_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08746_ _08745_/Y _08565_/X _06188_/X _08742_/X vssd1 vssd1 vccd1 vccd1 _12684_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _11845_/X _08670_/X _12711_/Q _08671_/X vssd1 vssd1 vccd1 vccd1 _12711_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _12951_/Q _12950_/Q _07650_/D vssd1 vssd1 vccd1 vccd1 _07658_/B sky130_fd_sc_hd__or3_4
XPHY_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07559_ _07558_/X _07552_/X _12991_/Q _07553_/X _07556_/X vssd1 vssd1 vccd1 vccd1
+ _12991_/D sky130_fd_sc_hd__a221o_1
XFILLER_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10570_ _10570_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _10570_/Y sky130_fd_sc_hd__nor2_1
XFILLER_166_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ _09229_/A vssd1 vssd1 vccd1 vccd1 _11675_/S sky130_fd_sc_hd__buf_4
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12240_ _12239_/X _12640_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12240_/X sky130_fd_sc_hd__mux2_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12171_ _11134_/X _10778_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _12171_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11122_ _10730_/X _11071_/A _06362_/X _11058_/A _12087_/X vssd1 vssd1 vccd1 vccd1
+ _11122_/X sky130_fd_sc_hd__a221o_1
XFILLER_122_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11053_ _11041_/X _11037_/X _06392_/X _07020_/X _11038_/X vssd1 vssd1 vccd1 vccd1
+ _11053_/X sky130_fd_sc_hd__a221o_1
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10004_ _08770_/Y _10003_/X _06227_/Y _10000_/X _10001_/X vssd1 vssd1 vccd1 vccd1
+ _10004_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_153_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11955_ _09861_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11955_/X sky130_fd_sc_hd__mux2_1
X_10906_ _12528_/Q vssd1 vssd1 vccd1 vccd1 _10906_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11886_ _11046_/X _11042_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _11886_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10837_ _12518_/Q vssd1 vssd1 vccd1 vccd1 _10837_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10768_ _11100_/A vssd1 vssd1 vccd1 vccd1 _10768_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12507_ _12509_/CLK _12507_/D vssd1 vssd1 vccd1 vccd1 _12507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10699_ _10699_/A vssd1 vssd1 vccd1 vccd1 _10699_/X sky130_fd_sc_hd__buf_2
XFILLER_145_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12438_ _12442_/CLK _12438_/D vssd1 vssd1 vccd1 vccd1 _12438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput406 _11188_/LO vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput417 _11198_/LO vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput428 _11208_/LO vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput439 _12771_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__clkbuf_2
X_12369_ _12369_/CLK _12369_/D vssd1 vssd1 vccd1 vccd1 _12369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06930_ _12001_/X _11998_/X _06924_/X _06925_/X _06929_/X vssd1 vssd1 vccd1 vccd1
+ _06931_/A sky130_fd_sc_hd__o32a_1
XFILLER_132_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06861_ _11111_/A _06861_/B vssd1 vssd1 vccd1 vccd1 _06861_/X sky130_fd_sc_hd__or2_1
XFILLER_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08600_ _08606_/A vssd1 vssd1 vccd1 vccd1 _08600_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06792_ _13199_/Q vssd1 vssd1 vccd1 vccd1 _06792_/Y sky130_fd_sc_hd__inv_2
X_09580_ _09592_/A _09580_/B vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__or2_1
XFILLER_94_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08531_ _11034_/A vssd1 vssd1 vccd1 vccd1 _10701_/A sky130_fd_sc_hd__buf_2
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08462_ _13065_/Q _10380_/A _08461_/Y _10318_/A vssd1 vssd1 vccd1 vccd1 _08467_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07413_ _07474_/A vssd1 vssd1 vccd1 vccd1 _07475_/A sky130_fd_sc_hd__inv_2
X_08393_ _08405_/A vssd1 vssd1 vccd1 vccd1 _08393_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07344_ _11441_/X _07338_/X _13065_/Q _07339_/X vssd1 vssd1 vccd1 vccd1 _13065_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07275_ _11550_/X _07263_/X _13085_/Q _07264_/X vssd1 vssd1 vccd1 vccd1 _13085_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09014_ _09016_/A _09016_/B _11640_/X vssd1 vssd1 vccd1 vccd1 _12584_/D sky130_fd_sc_hd__and3_1
X_06226_ _06245_/A vssd1 vssd1 vccd1 vccd1 _06226_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06157_ _12748_/Q _12716_/Q _06155_/X _06156_/X vssd1 vssd1 vccd1 vccd1 _06157_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06088_ _12695_/Q vssd1 vssd1 vccd1 vccd1 _06088_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09916_ _09939_/B vssd1 vssd1 vccd1 vccd1 _09935_/B sky130_fd_sc_hd__buf_1
XFILLER_113_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09847_ _09847_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _09868_/A sky130_fd_sc_hd__or2_2
XFILLER_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09778_ _13238_/Q _09777_/A _09686_/A _09777_/Y vssd1 vssd1 vccd1 vccd1 _09779_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _08729_/A vssd1 vssd1 vccd1 vccd1 _08729_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _09184_/A _11739_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11740_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11389_/X _09185_/B _11675_/S vssd1 vssd1 vccd1 vccd1 _11671_/X sky130_fd_sc_hd__mux2_1
XPHY_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10622_ _12414_/D _10620_/Y _09399_/Y _10620_/A _10617_/Y vssd1 vssd1 vccd1 vccd1
+ _10622_/X sky130_fd_sc_hd__o221a_1
XPHY_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10553_ _11393_/X vssd1 vssd1 vccd1 vccd1 _10553_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13272_ _13276_/CLK _13272_/D _06257_/X vssd1 vssd1 vccd1 vccd1 _13272_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10484_ _10484_/A _10484_/B vssd1 vssd1 vccd1 vccd1 _10486_/A sky130_fd_sc_hd__nand2_1
XFILLER_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12223_ _06300_/Y _13157_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12154_ _10007_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12154_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11105_ _10767_/X _11075_/X _06383_/X _11083_/X _11084_/X vssd1 vssd1 vccd1 vccd1
+ _11105_/X sky130_fd_sc_hd__a221o_1
XFILLER_2_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12085_ _12084_/X _12447_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12085_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11036_ _11036_/A vssd1 vssd1 vccd1 vccd1 _11036_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12987_ _12987_/CLK _12987_/D vssd1 vssd1 vccd1 vccd1 _12987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11938_ _09613_/Y _12799_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11938_/X sky130_fd_sc_hd__mux2_2
XFILLER_73_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11869_ _10192_/Y _12811_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11869_/X sky130_fd_sc_hd__mux2_1
XPHY_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07060_ _07053_/X _07058_/X _06305_/X _13156_/Q _07059_/X vssd1 vssd1 vccd1 vccd1
+ _13156_/D sky130_fd_sc_hd__a32o_1
XFILLER_199_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06011_ _06011_/A vssd1 vssd1 vccd1 vccd1 _09434_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_161_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07962_ _12895_/Q _11484_/X _07962_/S vssd1 vssd1 vccd1 vccd1 _12895_/D sky130_fd_sc_hd__mux2_1
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09701_ _09701_/A vssd1 vssd1 vccd1 vccd1 _09701_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06913_ _06917_/A _06918_/B vssd1 vssd1 vccd1 vccd1 _06913_/X sky130_fd_sc_hd__or2_1
X_07893_ _07967_/S vssd1 vssd1 vccd1 vccd1 _07904_/S sky130_fd_sc_hd__buf_2
XFILLER_96_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09632_ _09632_/A _09632_/B _09582_/A vssd1 vssd1 vccd1 vccd1 _09632_/X sky130_fd_sc_hd__or3b_1
X_06844_ _13192_/Q vssd1 vssd1 vccd1 vccd1 _06844_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09563_ _09563_/A vssd1 vssd1 vccd1 vccd1 _09563_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06775_ _06770_/X _06771_/X _06762_/X _06754_/X _06774_/X vssd1 vssd1 vccd1 vccd1
+ _06775_/X sky130_fd_sc_hd__o221a_1
XFILLER_43_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08514_ _12945_/Q vssd1 vssd1 vccd1 vccd1 _08514_/X sky130_fd_sc_hd__clkbuf_2
X_09494_ _12863_/Q vssd1 vssd1 vccd1 vccd1 _09494_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08445_ _13045_/Q vssd1 vssd1 vccd1 vccd1 _08445_/Y sky130_fd_sc_hd__inv_2
XPHY_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08376_ _12797_/Q _08374_/X _07997_/X _08375_/X vssd1 vssd1 vccd1 vccd1 _12797_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07327_ _11448_/X _07321_/X _13072_/Q _07324_/X vssd1 vssd1 vccd1 vccd1 _13072_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07258_ _07266_/A vssd1 vssd1 vccd1 vccd1 _07258_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06209_ _06209_/A _06209_/B _06209_/C _06253_/A vssd1 vssd1 vccd1 vccd1 _06209_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_118_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07189_ _11517_/X _07176_/X _13116_/Q _07177_/X vssd1 vssd1 vccd1 vccd1 _13116_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12910_ _12166_/X _12910_/D _07925_/X vssd1 vssd1 vccd1 vccd1 _12910_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_24_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12841_ _12166_/A0 _12841_/D _08255_/X vssd1 vssd1 vccd1 vccd1 _12841_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12773_/CLK _12772_/D _08438_/X vssd1 vssd1 vccd1 vccd1 _12772_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_199_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _09179_/B _11722_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11723_/X sky130_fd_sc_hd__mux2_1
XPHY_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _10544_/Y _10543_/Y _11704_/S vssd1 vssd1 vccd1 vccd1 _12366_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10605_ _10607_/A _11400_/X vssd1 vssd1 vccd1 vccd1 _10605_/Y sky130_fd_sc_hd__nor2b_1
XPHY_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11585_ _10421_/Y input357/X _11592_/S vssd1 vssd1 vccd1 vccd1 _11585_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10536_ _10557_/B vssd1 vssd1 vccd1 vccd1 _10554_/B sky130_fd_sc_hd__buf_2
XFILLER_171_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13255_ _13256_/CLK _13255_/D _06349_/X vssd1 vssd1 vccd1 vccd1 _13255_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10467_ _10467_/A _10467_/B _10467_/C vssd1 vssd1 vccd1 vccd1 _10468_/A sky130_fd_sc_hd__or3_4
XFILLER_170_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12206_ _12205_/X _12623_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12206_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13186_ _13193_/CLK _13186_/D _06894_/X vssd1 vssd1 vccd1 vccd1 _13186_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_57_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12986_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10398_ _10397_/A _10397_/B _10372_/X _10399_/A vssd1 vssd1 vccd1 vccd1 _10398_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12137_ _06468_/A _10707_/Y _12766_/Q vssd1 vssd1 vccd1 vccd1 _12202_/S sky130_fd_sc_hd__mux2_8
XFILLER_111_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12068_ _12067_/X _12445_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12068_/X sky130_fd_sc_hd__mux2_1
X_11019_ _12358_/Q _11018_/C _12359_/Q vssd1 vssd1 vccd1 vccd1 _11020_/B sky130_fd_sc_hd__a21oi_1
XFILLER_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06560_ _06580_/A vssd1 vssd1 vccd1 vccd1 _06560_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_79_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06491_ _06491_/A _12764_/Q vssd1 vssd1 vccd1 vccd1 _11077_/A sky130_fd_sc_hd__or2b_2
XFILLER_127_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08230_ _13101_/Q _10454_/A _08229_/Y _12822_/Q vssd1 vssd1 vccd1 vccd1 _08232_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08161_ _13125_/Q _10433_/A _08159_/Y _08160_/X vssd1 vssd1 vccd1 vccd1 _08162_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07112_ _07176_/A vssd1 vssd1 vccd1 vccd1 _07160_/A sky130_fd_sc_hd__buf_4
XFILLER_118_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08092_ _08098_/A vssd1 vssd1 vccd1 vccd1 _08092_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_173_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07043_ _07037_/X _07040_/X _06271_/Y _13162_/Q _07042_/X vssd1 vssd1 vccd1 vccd1
+ _13162_/D sky130_fd_sc_hd__a32o_1
XFILLER_161_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08994_ _12596_/Q vssd1 vssd1 vccd1 vccd1 _11029_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07945_ _07945_/A vssd1 vssd1 vccd1 vccd1 _07945_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07876_ _13025_/Q _10362_/B _13028_/Q _10367_/A _07875_/X vssd1 vssd1 vccd1 vccd1
+ _07879_/C sky130_fd_sc_hd__o221a_1
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09615_ _06905_/Y _06909_/Y _06891_/Y _09600_/Y vssd1 vssd1 vccd1 vccd1 _09620_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06827_ _07026_/A vssd1 vssd1 vccd1 vccd1 _06863_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ _09546_/A vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06758_ _11996_/X _06756_/B _06756_/X vssd1 vssd1 vccd1 vccd1 _06758_/X sky130_fd_sc_hd__a21bo_1
XFILLER_71_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ _12614_/Q vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__inv_2
X_06689_ _06457_/X _06682_/X _06688_/Y _06480_/X _13209_/Q vssd1 vssd1 vccd1 vccd1
+ _13209_/D sky130_fd_sc_hd__a32o_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08428_ _12777_/Q _08417_/X _07558_/X _08418_/X vssd1 vssd1 vccd1 vccd1 _12777_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08359_ _08359_/A vssd1 vssd1 vccd1 vccd1 _08375_/A sky130_fd_sc_hd__inv_2
XFILLER_149_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ _10662_/X _09310_/X _11370_/S vssd1 vssd1 vccd1 vccd1 _11370_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10321_ _10318_/A _12893_/Q _10318_/Y _07822_/Y _10320_/X vssd1 vssd1 vccd1 vccd1
+ _10321_/X sky130_fd_sc_hd__o221a_1
XFILLER_125_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13040_ _12164_/X _13040_/D _07408_/X vssd1 vssd1 vccd1 vccd1 _13040_/Q sky130_fd_sc_hd__dfrtp_4
X_10252_ _12888_/Q vssd1 vssd1 vccd1 vccd1 _10252_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10183_ _12629_/Q vssd1 vssd1 vccd1 vccd1 _10183_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12824_ _12169_/X _12824_/D _08306_/X vssd1 vssd1 vccd1 vccd1 _12824_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12755_ _13241_/CLK _12755_/D _08533_/X vssd1 vssd1 vccd1 vccd1 _12755_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11706_ _11705_/X _10627_/C _11774_/S vssd1 vssd1 vccd1 vccd1 _12417_/D sky130_fd_sc_hd__mux2_1
XPHY_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12719_/CLK _12686_/D _08736_/X vssd1 vssd1 vccd1 vccd1 _12686_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11637_ _10507_/X _12990_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11637_/X sky130_fd_sc_hd__mux2_1
XPHY_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11568_ _12825_/Q _09180_/A _11569_/S vssd1 vssd1 vccd1 vccd1 _11568_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10519_ _12396_/D _12397_/D vssd1 vssd1 vccd1 vccd1 _10561_/A sky130_fd_sc_hd__or2_1
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11499_ _10365_/Y _09179_/A _11501_/S vssd1 vssd1 vccd1 vccd1 _11499_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13238_ _13254_/CLK _13238_/D _06412_/X vssd1 vssd1 vccd1 vccd1 _13238_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_171_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13169_ _13170_/CLK _13169_/D _07016_/X vssd1 vssd1 vccd1 vccd1 _13169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07730_ _12611_/Q vssd1 vssd1 vccd1 vccd1 _09546_/A sky130_fd_sc_hd__inv_2
XFILLER_133_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07661_ _07661_/A _12961_/Q _07661_/C _12960_/Q vssd1 vssd1 vccd1 vccd1 _07689_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_81_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09400_ _09335_/Y _12397_/D _09354_/Y _12400_/D vssd1 vssd1 vccd1 vccd1 _09400_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06612_ _11894_/X _11892_/X _11894_/X _11892_/X vssd1 vssd1 vccd1 vccd1 _06612_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07592_ _09271_/C vssd1 vssd1 vccd1 vccd1 _09268_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09331_ _09331_/A _09331_/B vssd1 vssd1 vccd1 vccd1 _10548_/A sky130_fd_sc_hd__or2_1
XFILLER_179_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06543_ _06541_/X _06542_/X _06541_/X _06542_/X vssd1 vssd1 vccd1 vccd1 _06543_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_178_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09262_ _09284_/A _09279_/B _09260_/X _07508_/Y _09261_/X vssd1 vssd1 vccd1 vccd1
+ _09262_/X sky130_fd_sc_hd__o32a_1
X_06474_ _11883_/X _10787_/A _06473_/X vssd1 vssd1 vccd1 vccd1 _06474_/X sky130_fd_sc_hd__o21a_1
X_08213_ _13099_/Q vssd1 vssd1 vccd1 vccd1 _08213_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09193_ _12492_/Q _09190_/X _09179_/C _09192_/X vssd1 vssd1 vccd1 vccd1 _12492_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08144_ _12832_/Q vssd1 vssd1 vccd1 vccd1 _10480_/A sky130_fd_sc_hd__inv_2
XFILLER_14_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08075_ _08085_/A vssd1 vssd1 vccd1 vccd1 _08075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07026_ _07026_/A vssd1 vssd1 vccd1 vccd1 _07046_/A sky130_fd_sc_hd__buf_2
XFILLER_143_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput306 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _07101_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_103_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput317 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 _07100_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_102_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08977_ _09002_/A _08977_/B vssd1 vssd1 vccd1 vccd1 _12604_/D sky130_fd_sc_hd__nor2_1
Xinput328 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _09267_/B sky130_fd_sc_hd__clkbuf_4
Xinput339 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 input339/X sky130_fd_sc_hd__buf_2
XFILLER_25_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_2_wb_clk_i _12844_/CLK vssd1 vssd1 vccd1 vccd1 _12840_/CLK sky130_fd_sc_hd__clkbuf_16
X_07928_ _12909_/Q _11498_/X _07932_/S vssd1 vssd1 vccd1 vccd1 _12909_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07859_ _13036_/Q _10390_/A _07816_/Y _12902_/Q vssd1 vssd1 vccd1 vccd1 _07859_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ _10890_/A _10869_/X _10890_/A _10869_/X vssd1 vssd1 vccd1 vccd1 _12334_/D
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09555_/A vssd1 vssd1 vccd1 vccd1 _09530_/B sky130_fd_sc_hd__inv_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _12540_/CLK _12540_/D vssd1 vssd1 vccd1 vccd1 _12540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12471_ _12471_/CLK _12471_/D vssd1 vssd1 vccd1 vccd1 _12471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11422_ _12897_/Q input355/X _11422_/S vssd1 vssd1 vccd1 vccd1 _11422_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11353_ _09459_/X _12990_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _12317_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _10299_/Y _10163_/A _10300_/Y _10165_/A _10303_/X vssd1 vssd1 vccd1 vccd1
+ _10304_/X sky130_fd_sc_hd__o221a_1
XFILLER_125_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11284_ vssd1 vssd1 vccd1 vccd1 _11284_/HI _11284_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13023_ _12164_/X _13023_/D _07456_/X vssd1 vssd1 vccd1 vccd1 _13023_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10235_ _12782_/Q vssd1 vssd1 vccd1 vccd1 _10235_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10166_ _10166_/A vssd1 vssd1 vccd1 vccd1 _10166_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10097_ _10095_/Y _10018_/X _10096_/Y _10020_/X vssd1 vssd1 vccd1 vccd1 _10107_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12807_ _12169_/X _12807_/D _08346_/X vssd1 vssd1 vccd1 vccd1 _12807_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10999_ _12354_/Q vssd1 vssd1 vccd1 vccd1 _11014_/A sky130_fd_sc_hd__inv_2
XFILLER_37_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12738_ _12743_/CLK _12738_/D _08604_/X vssd1 vssd1 vccd1 vccd1 _12738_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_128_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12669_ _12683_/CLK _12669_/D _08796_/X vssd1 vssd1 vccd1 vccd1 _12669_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06190_ _06214_/A vssd1 vssd1 vccd1 vccd1 _06190_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_72_wb_clk_i _12960_/CLK vssd1 vssd1 vccd1 vccd1 _12957_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08900_ _08963_/A vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__clkbuf_2
X_09880_ _09880_/A _09880_/B vssd1 vssd1 vccd1 vccd1 _09881_/B sky130_fd_sc_hd__or2_1
XFILLER_135_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08831_ _08814_/A _08781_/A _06342_/Y _12656_/Q _08567_/A vssd1 vssd1 vccd1 vccd1
+ _12656_/D sky130_fd_sc_hd__a32o_1
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08762_ _08769_/A vssd1 vssd1 vccd1 vccd1 _08762_/X sky130_fd_sc_hd__clkbuf_1
X_07713_ _12954_/Q _07707_/X _12953_/Q _07705_/X _07703_/X vssd1 vssd1 vccd1 vccd1
+ _12954_/D sky130_fd_sc_hd__o221a_1
XFILLER_54_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08693_ _08699_/A vssd1 vssd1 vccd1 vccd1 _08693_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07644_ _07660_/D _07650_/D vssd1 vssd1 vccd1 vccd1 _07689_/B sky130_fd_sc_hd__or2_2
XPHY_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07575_ _07575_/A vssd1 vssd1 vccd1 vccd1 _07575_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09314_ _09314_/A vssd1 vssd1 vccd1 vccd1 _12139_/S sky130_fd_sc_hd__inv_4
X_06526_ _06886_/A vssd1 vssd1 vccd1 vccd1 _06526_/X sky130_fd_sc_hd__buf_2
XFILLER_181_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09245_ _10528_/A _09245_/B _10529_/B _10528_/B vssd1 vssd1 vccd1 vccd1 _09246_/A
+ sky130_fd_sc_hd__or4b_4
X_06457_ _06887_/A vssd1 vssd1 vccd1 vccd1 _06457_/X sky130_fd_sc_hd__buf_4
XFILLER_178_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09176_ _11029_/A _09175_/B _12595_/Q _12493_/Q _09175_/Y vssd1 vssd1 vccd1 vccd1
+ _12493_/D sky130_fd_sc_hd__a32o_1
X_06388_ _06391_/A vssd1 vssd1 vccd1 vccd1 _06388_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08127_ _13135_/Q vssd1 vssd1 vccd1 vccd1 _08127_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08058_ _12863_/Q _08040_/A _07304_/X _08041_/A vssd1 vssd1 vccd1 vccd1 _12863_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07009_ _06886_/X _07008_/X _06887_/X _13172_/Q vssd1 vssd1 vccd1 vccd1 _13172_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_89_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10020_ _10163_/A vssd1 vssd1 vccd1 vccd1 _10020_/X sky130_fd_sc_hd__clkbuf_2
Xinput103 la_data_in[42] vssd1 vssd1 vccd1 vccd1 input103/X sky130_fd_sc_hd__buf_1
XFILLER_103_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput114 la_data_in[52] vssd1 vssd1 vccd1 vccd1 input114/X sky130_fd_sc_hd__buf_1
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput125 la_data_in[62] vssd1 vssd1 vccd1 vccd1 input125/X sky130_fd_sc_hd__buf_1
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput136 la_data_in[72] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_hd__buf_1
Xinput147 la_data_in[82] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_hd__buf_1
XFILLER_130_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput158 la_data_in[92] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_hd__buf_1
Xinput169 la_oenb[101] vssd1 vssd1 vccd1 vccd1 input169/X sky130_fd_sc_hd__buf_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11971_ _12973_/Q _12925_/Q _12602_/Q vssd1 vssd1 vccd1 vccd1 _11971_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10922_ _10911_/Y _10912_/Y _10906_/Y _10907_/Y vssd1 vssd1 vccd1 vccd1 _10922_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10853_ _10851_/X _10852_/X _10851_/X _10852_/X vssd1 vssd1 vccd1 vccd1 _12332_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_201_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _10736_/X _10768_/X _06365_/X _10769_/X _10770_/X vssd1 vssd1 vccd1 vccd1
+ _10784_/X sky130_fd_sc_hd__a221o_1
XFILLER_188_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12523_ _12802_/CLK _12523_/D vssd1 vssd1 vccd1 vccd1 _12523_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12454_ _12455_/CLK _12454_/D vssd1 vssd1 vccd1 vccd1 _12454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11405_ _10616_/Y _12411_/D _11889_/S vssd1 vssd1 vccd1 vccd1 _11405_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ _12472_/CLK _12385_/D vssd1 vssd1 vccd1 vccd1 _12407_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_138_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11336_ vssd1 vssd1 vccd1 vccd1 _11336_/HI _11336_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11267_ vssd1 vssd1 vccd1 vccd1 _11267_/HI _11267_/LO sky130_fd_sc_hd__conb_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13006_ _13008_/CLK _13006_/D vssd1 vssd1 vccd1 vccd1 _13006_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10218_ _12781_/Q vssd1 vssd1 vccd1 vccd1 _10218_/Y sky130_fd_sc_hd__inv_2
X_11198_ vssd1 vssd1 vccd1 vccd1 _11198_/HI _11198_/LO sky130_fd_sc_hd__conb_1
XFILLER_95_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10149_ _09906_/Y _10134_/X _10138_/X _10148_/X vssd1 vssd1 vccd1 vccd1 _10149_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07360_ _07360_/A vssd1 vssd1 vccd1 vccd1 _07360_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06311_ _06311_/A vssd1 vssd1 vccd1 vccd1 _06311_/Y sky130_fd_sc_hd__clkinv_4
X_07291_ _13080_/Q _07285_/X _07290_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _13080_/D
+ sky130_fd_sc_hd__a22o_1
X_09030_ _09030_/A vssd1 vssd1 vccd1 vccd1 _09030_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06242_ _06053_/Y _06054_/Y _06241_/Y _06196_/X vssd1 vssd1 vccd1 vccd1 _06242_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_191_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06173_ _06079_/Y _06182_/B _06140_/X vssd1 vssd1 vccd1 vccd1 _06173_/X sky130_fd_sc_hd__o21a_1
XFILLER_172_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09932_ _12890_/Q _09935_/B vssd1 vssd1 vccd1 vccd1 _09932_/X sky130_fd_sc_hd__or2_1
XFILLER_104_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09863_ _13236_/Q _13235_/Q _09862_/Y _06441_/Y vssd1 vssd1 vccd1 vccd1 _09864_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_97_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08814_ _08814_/A vssd1 vssd1 vccd1 vccd1 _08814_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09794_ _09794_/A vssd1 vssd1 vccd1 vccd1 _09794_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08745_ _12684_/Q vssd1 vssd1 vccd1 vccd1 _08745_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08676_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08676_/X sky130_fd_sc_hd__clkbuf_1
XPHY_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07664_/A _07660_/C vssd1 vssd1 vccd1 vccd1 _07650_/D sky130_fd_sc_hd__or2_1
XPHY_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ _09185_/B vssd1 vssd1 vccd1 vccd1 _07558_/X sky130_fd_sc_hd__buf_4
XFILLER_167_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06509_ _12160_/X vssd1 vssd1 vccd1 vccd1 _06509_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07489_ _07489_/A vssd1 vssd1 vccd1 vccd1 _07489_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09228_ _09228_/A _09228_/B _09228_/C _10558_/B vssd1 vssd1 vccd1 vccd1 _09229_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_166_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09159_ _11632_/X _09154_/X _12507_/Q _09156_/X vssd1 vssd1 vccd1 vccd1 _12507_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12170_ _11140_/X _11139_/Y _12193_/S vssd1 vssd1 vccd1 vccd1 _12170_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11121_ _10693_/X _10737_/X _06407_/X _10738_/X _10739_/X vssd1 vssd1 vccd1 vccd1
+ _11121_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11052_ _06386_/X _11045_/X _11032_/X _10773_/X _11034_/X vssd1 vssd1 vccd1 vccd1
+ _11052_/X sky130_fd_sc_hd__a32o_1
XFILLER_67_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10003_ _10003_/A vssd1 vssd1 vccd1 vccd1 _10003_/X sky130_fd_sc_hd__buf_2
XFILLER_49_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11954_ _09855_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11954_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10905_ _10903_/A _10904_/A _10921_/B _10904_/Y vssd1 vssd1 vccd1 vccd1 _12339_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11885_ _10743_/X _10791_/X _12193_/S vssd1 vssd1 vccd1 vccd1 _11885_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10836_ _10827_/A _10831_/Y _10828_/A _10835_/X vssd1 vssd1 vccd1 vccd1 _10836_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_199_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10767_ _10767_/A vssd1 vssd1 vccd1 vccd1 _10767_/X sky130_fd_sc_hd__buf_2
XFILLER_201_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12506_ _12509_/CLK _12506_/D vssd1 vssd1 vccd1 vccd1 _12506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ _13242_/Q vssd1 vssd1 vccd1 vccd1 _10699_/A sky130_fd_sc_hd__inv_2
XFILLER_195_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12437_ _12441_/CLK _12437_/D vssd1 vssd1 vccd1 vccd1 _12437_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_201_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput407 _11189_/LO vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__clkbuf_2
Xoutput418 _11199_/LO vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__clkbuf_2
X_12368_ _12369_/CLK _12368_/D vssd1 vssd1 vccd1 vccd1 _12368_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput429 _11209_/LO vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11319_ vssd1 vssd1 vccd1 vccd1 _11319_/HI _11319_/LO sky130_fd_sc_hd__conb_1
X_12299_ _12977_/CLK _12299_/D vssd1 vssd1 vccd1 vccd1 _12299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06860_ _06860_/A vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06791_ _12016_/X _12012_/X _06785_/X _06786_/X _06790_/X vssd1 vssd1 vccd1 vccd1
+ _06791_/X sky130_fd_sc_hd__o32a_2
XFILLER_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08530_ _08533_/A vssd1 vssd1 vccd1 vccd1 _08530_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08461_ _13043_/Q vssd1 vssd1 vccd1 vccd1 _08461_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07412_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07412_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08392_ _12790_/Q _08374_/A _07304_/X _08375_/A vssd1 vssd1 vccd1 vccd1 _12790_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07343_ _07345_/A vssd1 vssd1 vccd1 vccd1 _07343_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07274_ _07280_/A vssd1 vssd1 vccd1 vccd1 _07274_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09013_ _09016_/A _09016_/B _11641_/X vssd1 vssd1 vccd1 vccd1 _12585_/D sky130_fd_sc_hd__and3_1
XFILLER_136_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06225_ _06222_/Y _06216_/X _06217_/X _06224_/X vssd1 vssd1 vccd1 vccd1 _13279_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06156_ _12748_/Q _12716_/Q _12747_/Q _12715_/Q vssd1 vssd1 vccd1 vccd1 _06156_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06087_ _12727_/Q vssd1 vssd1 vccd1 vccd1 _06087_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09915_ _09949_/A vssd1 vssd1 vccd1 vccd1 _09915_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09846_ _06462_/Y _09845_/X _06462_/Y _09845_/X vssd1 vssd1 vccd1 vccd1 _09866_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_101_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09777_ _09777_/A vssd1 vssd1 vccd1 vccd1 _09777_/Y sky130_fd_sc_hd__inv_2
X_06989_ _11882_/X vssd1 vssd1 vccd1 vccd1 _06989_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _11824_/X _08715_/X _12690_/Q _08716_/X vssd1 vssd1 vccd1 vccd1 _12690_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08659_ _08669_/A vssd1 vssd1 vccd1 vccd1 _08659_/X sky130_fd_sc_hd__clkbuf_1
XPHY_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11669_/X _11392_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12377_/D sky130_fd_sc_hd__mux2_1
XPHY_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _10619_/A _10619_/B _10620_/Y _10617_/A vssd1 vssd1 vccd1 vccd1 _10621_/Y
+ sky130_fd_sc_hd__a211oi_2
XPHY_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10552_ _12369_/Q _10548_/Y _09333_/B vssd1 vssd1 vccd1 vccd1 _10552_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_183_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13271_ _13276_/CLK _13271_/D _06262_/X vssd1 vssd1 vccd1 vccd1 _13271_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10483_ _10482_/A _10482_/B _10474_/A _10484_/B vssd1 vssd1 vccd1 vccd1 _10483_/Y
+ sky130_fd_sc_hd__a211oi_2
Xclkbuf_leaf_129_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13256_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12222_ _12221_/X _12631_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__mux2_2
XFILLER_154_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12153_ _10006_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12153_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _10758_/X _11054_/A _06376_/X _11055_/A _11899_/X vssd1 vssd1 vccd1 vccd1
+ _11104_/X sky130_fd_sc_hd__a221o_1
XFILLER_151_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12084_ _12447_/Q _12083_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11035_ _06397_/X _10691_/A _11032_/X _11033_/X _11034_/X vssd1 vssd1 vccd1 vccd1
+ _11035_/X sky130_fd_sc_hd__a32o_1
XFILLER_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12986_ _12986_/CLK _12986_/D vssd1 vssd1 vccd1 vccd1 _12986_/Q sky130_fd_sc_hd__dfxtp_1
X_11937_ _09597_/X _12798_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11937_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11868_ _10173_/Y _12319_/Q _12312_/Q vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__mux2_2
XFILLER_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10819_ _10814_/Y _10815_/Y _10821_/C _10821_/A vssd1 vssd1 vccd1 vccd1 _10819_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11799_ _12065_/X _12484_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11799_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06010_ _09986_/D _09981_/C _09433_/A _06011_/A vssd1 vssd1 vccd1 vccd1 _06017_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_173_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07961_ _07961_/A vssd1 vssd1 vccd1 vccd1 _07961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09700_ _09700_/A _09700_/B vssd1 vssd1 vccd1 vccd1 _09700_/X sky130_fd_sc_hd__or2_1
X_06912_ _06910_/X _06911_/X _06910_/X _06911_/X vssd1 vssd1 vccd1 vccd1 _06918_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_136_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07892_ _07951_/A vssd1 vssd1 vccd1 vccd1 _07967_/S sky130_fd_sc_hd__buf_4
XFILLER_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09631_ _09614_/Y _09630_/A _09621_/Y vssd1 vssd1 vccd1 vccd1 _09675_/A sky130_fd_sc_hd__o21ai_1
X_06843_ _06863_/A vssd1 vssd1 vccd1 vccd1 _06843_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09562_ _13180_/Q _13179_/Q _09578_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09563_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_167_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06774_ _06778_/A _06778_/B vssd1 vssd1 vccd1 vccd1 _06774_/X sky130_fd_sc_hd__or2_1
XFILLER_24_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08513_ _08518_/A vssd1 vssd1 vccd1 vccd1 _08513_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09493_ _09490_/A _09490_/B _09492_/X vssd1 vssd1 vccd1 vccd1 _09493_/Y sky130_fd_sc_hd__o21ai_1
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08444_ _08440_/Y _12897_/Q _13046_/Q _10328_/A _08443_/X vssd1 vssd1 vccd1 vccd1
+ _08457_/A sky130_fd_sc_hd__a221o_1
XPHY_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ _08375_/A vssd1 vssd1 vccd1 vccd1 _08375_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07326_ _07330_/A vssd1 vssd1 vccd1 vccd1 _07326_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07257_ _11557_/X _07248_/X _13092_/Q _07249_/X vssd1 vssd1 vccd1 vccd1 _13092_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06208_ _06182_/A _06182_/B _06181_/X _06173_/X vssd1 vssd1 vccd1 vccd1 _06253_/A
+ sky130_fd_sc_hd__o31a_1
X_07188_ _07206_/A vssd1 vssd1 vccd1 vccd1 _07188_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06139_ _06209_/A _06136_/Y _06138_/Y vssd1 vssd1 vccd1 vccd1 _06197_/A sky130_fd_sc_hd__o21a_1
XFILLER_155_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09829_ _09829_/A _09868_/C vssd1 vssd1 vccd1 vccd1 _09829_/X sky130_fd_sc_hd__or2_1
XFILLER_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12840_ _12840_/CLK _12840_/D _08257_/X vssd1 vssd1 vccd1 vccd1 _12840_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_100_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12771_ _12169_/A0 _12771_/D vssd1 vssd1 vccd1 vccd1 _12771_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11915_/X _12485_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11722_/X sky130_fd_sc_hd__mux2_1
XPHY_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _10540_/Y _10539_/Y _11704_/S vssd1 vssd1 vccd1 vccd1 _12365_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10604_ _12409_/D _10602_/Y _10603_/X vssd1 vssd1 vccd1 vccd1 _10604_/X sky130_fd_sc_hd__o21a_1
XPHY_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11584_ _10419_/X _09185_/B _11592_/S vssd1 vssd1 vccd1 vccd1 _11584_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10535_ _10535_/A vssd1 vssd1 vccd1 vccd1 _10557_/B sky130_fd_sc_hd__inv_2
XPHY_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13254_ _13254_/CLK _13254_/D _06353_/X vssd1 vssd1 vccd1 vccd1 _13254_/Q sky130_fd_sc_hd__dfrtp_2
X_10466_ _10467_/B _10467_/C _12826_/Q _10464_/A _10437_/X vssd1 vssd1 vccd1 vccd1
+ _10466_/X sky130_fd_sc_hd__o221a_1
XFILLER_171_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12205_ _06346_/Y _13148_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12205_/X sky130_fd_sc_hd__mux2_1
X_13185_ _13190_/CLK _13185_/D _06908_/X vssd1 vssd1 vccd1 vccd1 _13185_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10397_ _10397_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10399_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12136_ _12135_/X _12435_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12136_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12067_ _12445_/Q _12066_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _12067_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_97_wb_clk_i _13235_/CLK vssd1 vssd1 vccd1 vccd1 _13190_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11018_ _12358_/Q _12359_/Q _11018_/C vssd1 vssd1 vccd1 vccd1 _11021_/B sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_26_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12480_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12969_ _12984_/CLK _12969_/D vssd1 vssd1 vccd1 vccd1 _12969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06490_ _12763_/Q _12762_/Q vssd1 vssd1 vccd1 vccd1 _06491_/A sky130_fd_sc_hd__and2_1
XFILLER_127_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08160_ _12812_/Q vssd1 vssd1 vccd1 vccd1 _08160_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07111_ hold1/X _11546_/S vssd1 vssd1 vccd1 vccd1 _07176_/A sky130_fd_sc_hd__or2_1
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08091_ _12851_/Q _08082_/X _08005_/X _08083_/X vssd1 vssd1 vccd1 vccd1 _12851_/D
+ sky130_fd_sc_hd__a22o_1
X_07042_ _07042_/A vssd1 vssd1 vccd1 vccd1 _07042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08993_ _12599_/Q _12598_/Q _09019_/A _08992_/Y vssd1 vssd1 vccd1 vccd1 _12599_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07944_ _12902_/Q _11491_/X _07946_/S vssd1 vssd1 vccd1 vccd1 _12902_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07875_ _13038_/Q _10395_/A _13022_/Q _10352_/A vssd1 vssd1 vccd1 vccd1 _07875_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_56_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09614_ _09614_/A vssd1 vssd1 vccd1 vccd1 _09614_/Y sky130_fd_sc_hd__inv_2
X_06826_ _07477_/A vssd1 vssd1 vccd1 vccd1 _07026_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09545_ _09939_/B vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__buf_2
X_06757_ _12002_/X _11999_/X _06756_/X vssd1 vssd1 vccd1 vccd1 _06757_/X sky130_fd_sc_hd__o21a_1
XFILLER_36_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09476_ _12861_/Q vssd1 vssd1 vccd1 vccd1 _09476_/Y sky130_fd_sc_hd__inv_2
X_06688_ _12199_/X _06688_/B vssd1 vssd1 vccd1 vccd1 _06688_/Y sky130_fd_sc_hd__nand2_1
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08427_ _08433_/A vssd1 vssd1 vccd1 vccd1 _08427_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_197_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08358_ _08374_/A vssd1 vssd1 vccd1 vccd1 _08358_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07309_ _09226_/B vssd1 vssd1 vccd1 vccd1 _07309_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_165_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08289_ _08296_/A vssd1 vssd1 vccd1 vccd1 _08289_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10320_ _10372_/A vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__buf_2
XFILLER_166_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10251_ _12783_/Q vssd1 vssd1 vccd1 vccd1 _10251_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10182_ _12884_/Q vssd1 vssd1 vccd1 vccd1 _10182_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput590 _12562_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12823_ _12169_/X _12823_/D _08308_/X vssd1 vssd1 vccd1 vccd1 _12823_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_27_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12942_/CLK _12754_/D _08539_/X vssd1 vssd1 vccd1 vccd1 _12754_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _10627_/C _10627_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11705_/X sky130_fd_sc_hd__mux2_1
XPHY_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12685_/CLK _12685_/D _08738_/X vssd1 vssd1 vccd1 vccd1 _12685_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_187_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_144_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12871_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11636_ _10506_/X _12989_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11636_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11567_ _12824_/Q _09180_/B _11569_/S vssd1 vssd1 vccd1 vccd1 _11567_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10518_ _12592_/Q _07766_/B _11648_/S vssd1 vssd1 vccd1 vccd1 _10518_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11498_ _10361_/X _09179_/B _11501_/S vssd1 vssd1 vccd1 vccd1 _11498_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13237_ _13237_/CLK _13237_/D _06417_/X vssd1 vssd1 vccd1 vccd1 _13237_/Q sky130_fd_sc_hd__dfrtp_1
X_10449_ _10455_/A _10449_/B _10455_/D vssd1 vssd1 vccd1 vccd1 _10450_/A sky130_fd_sc_hd__or3_4
XFILLER_170_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13168_ _13177_/CLK _13168_/D _07018_/X vssd1 vssd1 vccd1 vccd1 _13168_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12119_ _12118_/X _12436_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12119_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13099_ _12167_/X _13099_/D _07239_/X vssd1 vssd1 vccd1 vccd1 _13099_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07660_ _12959_/Q _12958_/Q _07660_/C _07660_/D vssd1 vssd1 vccd1 vccd1 _07661_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06611_ _11893_/X _11898_/X _06609_/X vssd1 vssd1 vccd1 vccd1 _06611_/X sky130_fd_sc_hd__a21bo_1
X_07591_ _09276_/C vssd1 vssd1 vccd1 vccd1 _09271_/C sky130_fd_sc_hd__inv_2
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _09330_/A _10541_/A vssd1 vssd1 vccd1 vccd1 _09331_/B sky130_fd_sc_hd__or2_1
X_06542_ _12176_/X _12175_/X _12176_/X _12175_/X vssd1 vssd1 vccd1 vccd1 _06542_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_179_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09261_ _09279_/A _09279_/D _13008_/Q _09276_/C vssd1 vssd1 vccd1 vccd1 _09261_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_179_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06473_ _11885_/X _06479_/B vssd1 vssd1 vccd1 vccd1 _06473_/X sky130_fd_sc_hd__or2_1
X_08212_ _08210_/Y _08160_/X _13082_/Q _08176_/Y _08211_/X vssd1 vssd1 vccd1 vccd1
+ _08222_/A sky130_fd_sc_hd__a221o_1
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09192_ _09216_/A vssd1 vssd1 vccd1 vccd1 _09192_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08143_ _13137_/Q _10467_/A _08141_/Y _10405_/A vssd1 vssd1 vccd1 vccd1 _08151_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08074_ _12858_/Q _08066_/X _07983_/X _08068_/X vssd1 vssd1 vccd1 vccd1 _12858_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07025_ _06663_/X _12183_/X _06415_/B _13166_/Q vssd1 vssd1 vccd1 vccd1 _13166_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_115_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput307 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _07515_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput318 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _11964_/S sky130_fd_sc_hd__buf_4
XFILLER_76_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08976_ _09002_/A _08976_/B vssd1 vssd1 vccd1 vccd1 _12605_/D sky130_fd_sc_hd__nor2_1
Xinput329 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 input329/X sky130_fd_sc_hd__clkbuf_2
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07927_ _07931_/A vssd1 vssd1 vccd1 vccd1 _07927_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07858_ _07858_/A _07858_/B _07858_/C _07857_/X vssd1 vssd1 vccd1 vccd1 _07867_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06809_ _11881_/X _06807_/Y _06808_/Y _11880_/X vssd1 vssd1 vccd1 vccd1 _06861_/B
+ sky130_fd_sc_hd__o22a_1
X_07789_ _07568_/X _07780_/A _12926_/Q _07781_/A _07522_/A vssd1 vssd1 vccd1 vccd1
+ _12926_/D sky130_fd_sc_hd__a221o_1
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09528_ _09528_/A _09528_/B vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__or2_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _13005_/Q _09442_/X _09457_/X _09458_/X vssd1 vssd1 vccd1 vccd1 _09459_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_52_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12470_ _12471_/CLK _12470_/D vssd1 vssd1 vccd1 vccd1 _12470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11421_ _12896_/Q _09186_/B _11422_/S vssd1 vssd1 vccd1 vccd1 _11421_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11352_ _09456_/X _12989_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _12316_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10303_ _10301_/Y _10166_/A _10302_/Y _10168_/A vssd1 vssd1 vccd1 vccd1 _10303_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11283_ vssd1 vssd1 vccd1 vccd1 _11283_/HI _11283_/LO sky130_fd_sc_hd__conb_1
XFILLER_106_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _12164_/X _13022_/D _07458_/X vssd1 vssd1 vccd1 vccd1 _13022_/Q sky130_fd_sc_hd__dfrtp_2
X_10234_ _10232_/Y _10032_/X _10233_/Y _10137_/X vssd1 vssd1 vccd1 vccd1 _10234_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10165_ _10165_/A vssd1 vssd1 vccd1 vccd1 _10165_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10096_ _12880_/Q vssd1 vssd1 vccd1 vccd1 _10096_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12806_ _12169_/X _12806_/D _08348_/X vssd1 vssd1 vccd1 vccd1 _12806_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10998_ _10995_/Y _10997_/A _11000_/D _10997_/Y vssd1 vssd1 vccd1 vccd1 _12353_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12737_ _12737_/CLK _12737_/D _08606_/X vssd1 vssd1 vccd1 vccd1 _12737_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_70_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12668_ _12683_/CLK _12668_/D _08800_/X vssd1 vssd1 vccd1 vccd1 _12668_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11619_ _10489_/Y _12986_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11619_/X sky130_fd_sc_hd__mux2_1
X_12599_ _12937_/CLK _12599_/D vssd1 vssd1 vccd1 vccd1 _12599_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_41_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13008_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08830_ _08836_/A vssd1 vssd1 vccd1 vccd1 _08830_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08761_ _08759_/Y _08760_/X _06212_/X _08742_/X vssd1 vssd1 vccd1 vccd1 _12680_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07712_ _12955_/Q _07707_/X _07698_/X _07711_/Y _07703_/X vssd1 vssd1 vccd1 vccd1
+ _12955_/D sky130_fd_sc_hd__o221a_1
X_08692_ _11839_/X _08685_/X _12705_/Q _08686_/X vssd1 vssd1 vccd1 vccd1 _12705_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07643_ _12962_/Q vssd1 vssd1 vccd1 vccd1 _07659_/A sky130_fd_sc_hd__inv_2
XFILLER_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07574_ _07574_/A vssd1 vssd1 vccd1 vccd1 _07574_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09313_ _12436_/Q _12435_/Q vssd1 vssd1 vccd1 vccd1 _09313_/X sky130_fd_sc_hd__or2_1
XFILLER_81_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06525_ _06580_/A vssd1 vssd1 vccd1 vccd1 _06525_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_181_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09244_ _09244_/A _09244_/B vssd1 vssd1 vccd1 vccd1 _10529_/B sky130_fd_sc_hd__nand2_2
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06456_ _06465_/A vssd1 vssd1 vccd1 vccd1 _06456_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ _11029_/A _09175_/B vssd1 vssd1 vccd1 vccd1 _09175_/Y sky130_fd_sc_hd__nand2_1
XFILLER_182_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06387_ _06382_/X _12218_/X _06375_/X _06386_/X vssd1 vssd1 vccd1 vccd1 _13246_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08126_ _12827_/Q vssd1 vssd1 vccd1 vccd1 _10467_/A sky130_fd_sc_hd__inv_2
XFILLER_147_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08057_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08057_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07008_ _11055_/A vssd1 vssd1 vccd1 vccd1 _07008_/X sky130_fd_sc_hd__buf_2
XFILLER_116_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput104 la_data_in[43] vssd1 vssd1 vccd1 vccd1 input104/X sky130_fd_sc_hd__buf_1
XFILLER_102_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput115 la_data_in[53] vssd1 vssd1 vccd1 vccd1 input115/X sky130_fd_sc_hd__buf_1
XFILLER_103_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput126 la_data_in[63] vssd1 vssd1 vccd1 vccd1 input126/X sky130_fd_sc_hd__buf_1
XFILLER_5_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput137 la_data_in[73] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_hd__buf_1
XFILLER_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput148 la_data_in[83] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_hd__buf_1
Xinput159 la_data_in[93] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_hd__buf_1
X_08959_ _08962_/A vssd1 vssd1 vccd1 vccd1 _08959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11970_ _07737_/X _09259_/Y _12607_/Q vssd1 vssd1 vccd1 vccd1 _11970_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10921_ _10921_/A _10921_/B _10921_/C _10908_/X vssd1 vssd1 vccd1 vccd1 _10944_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_99_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10852_ _12519_/Q _12331_/Q _10843_/Y _10846_/Y vssd1 vssd1 vccd1 vccd1 _10852_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10783_ _10730_/X _10768_/X _06362_/X _10769_/X _10770_/X vssd1 vssd1 vccd1 vccd1
+ _10783_/X sky130_fd_sc_hd__a221o_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12522_ _12801_/CLK _12522_/D vssd1 vssd1 vccd1 vccd1 _12522_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12453_ _12458_/CLK _12453_/D vssd1 vssd1 vccd1 vccd1 _12453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11404_ _10598_/Y _12407_/D _11404_/S vssd1 vssd1 vccd1 vccd1 _11404_/X sky130_fd_sc_hd__mux2_1
X_12384_ _12472_/CLK _12384_/D vssd1 vssd1 vccd1 vccd1 _12406_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11335_ vssd1 vssd1 vccd1 vccd1 _11335_/HI _11335_/LO sky130_fd_sc_hd__conb_1
XFILLER_67_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11266_ vssd1 vssd1 vccd1 vccd1 _11266_/HI _11266_/LO sky130_fd_sc_hd__conb_1
X_13005_ _13008_/CLK _13005_/D vssd1 vssd1 vccd1 vccd1 _13005_/Q sky130_fd_sc_hd__dfxtp_2
X_10217_ _10215_/Y _10000_/A _10216_/Y _10137_/X vssd1 vssd1 vccd1 vccd1 _10217_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11197_ vssd1 vssd1 vccd1 vccd1 _11197_/HI _11197_/LO sky130_fd_sc_hd__conb_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10148_ _10139_/Y _10140_/X _09532_/Y _10141_/X _10147_/X vssd1 vssd1 vccd1 vccd1
+ _10148_/X sky130_fd_sc_hd__o221a_1
XFILLER_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10079_ _12640_/Q vssd1 vssd1 vccd1 vccd1 _10079_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06310_ _06103_/A _06309_/X _06103_/A _06309_/X vssd1 vssd1 vccd1 vccd1 _06311_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_31_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07290_ _09185_/A vssd1 vssd1 vccd1 vccd1 _07290_/X sky130_fd_sc_hd__buf_2
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06241_ _06241_/A vssd1 vssd1 vccd1 vccd1 _06241_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06172_ _06172_/A _06172_/B vssd1 vssd1 vccd1 vccd1 _06209_/C sky130_fd_sc_hd__or2_1
XFILLER_116_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09931_ _12667_/Q vssd1 vssd1 vccd1 vccd1 _09931_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09862_ _13236_/Q vssd1 vssd1 vccd1 vccd1 _09862_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08813_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08813_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09793_ _09782_/A _09782_/B _09785_/X vssd1 vssd1 vccd1 vccd1 _09794_/A sky130_fd_sc_hd__o21ai_1
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08744_ _08747_/A vssd1 vssd1 vccd1 vccd1 _08744_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08675_ _11846_/X _08670_/X _12712_/Q _08671_/X vssd1 vssd1 vccd1 vccd1 _12712_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _12955_/Q _12954_/Q _12957_/Q _12956_/Q vssd1 vssd1 vccd1 vccd1 _07660_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07557_ _07536_/X _07552_/X _12992_/Q _07553_/X _07556_/X vssd1 vssd1 vccd1 vccd1
+ _12992_/D sky130_fd_sc_hd__a221o_1
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06508_ _13227_/Q vssd1 vssd1 vccd1 vccd1 _06508_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07488_ _11452_/X _07474_/X _13011_/Q _07475_/X vssd1 vssd1 vccd1 vccd1 _13011_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09227_ _09227_/A _09227_/B _07568_/A _07562_/A vssd1 vssd1 vccd1 vccd1 _10558_/B
+ sky130_fd_sc_hd__or4bb_4
X_06439_ _12621_/Q vssd1 vssd1 vccd1 vccd1 _06658_/A sky130_fd_sc_hd__buf_4
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09158_ _11633_/X _09154_/X _12508_/Q _09156_/X vssd1 vssd1 vccd1 vccd1 _12508_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08109_ _13116_/Q vssd1 vssd1 vccd1 vccd1 _08109_/Y sky130_fd_sc_hd__inv_2
X_09089_ _09115_/A vssd1 vssd1 vccd1 vccd1 _09089_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11120_ _10699_/A _10788_/X _13242_/Q _11111_/X _11112_/X vssd1 vssd1 vccd1 vccd1
+ _11120_/X sky130_fd_sc_hd__a221o_1
XFILLER_190_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11051_ _11051_/A vssd1 vssd1 vccd1 vccd1 _11051_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10002_ _08774_/Y _09993_/X _06231_/Y _10000_/X _10001_/X vssd1 vssd1 vccd1 vccd1
+ _10002_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11953_ _09843_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11953_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10904_ _10904_/A vssd1 vssd1 vccd1 vccd1 _10904_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11884_ _11044_/X _11040_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _11884_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ _10827_/A _10831_/Y _10828_/B _10834_/X vssd1 vssd1 vccd1 vccd1 _10835_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_198_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10766_ _13247_/Q vssd1 vssd1 vccd1 vccd1 _10767_/A sky130_fd_sc_hd__inv_2
XFILLER_185_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12505_ _13244_/CLK _12505_/D vssd1 vssd1 vccd1 vccd1 _12505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10697_ _06404_/X _10691_/A _10691_/B _10696_/X _10701_/A vssd1 vssd1 vccd1 vccd1
+ _10697_/X sky130_fd_sc_hd__a32o_1
XFILLER_186_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12436_ _12441_/CLK _12436_/D vssd1 vssd1 vccd1 vccd1 _12436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput408 _11190_/LO vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_153_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput419 _11200_/LO vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__clkbuf_2
X_12367_ _12369_/CLK _12367_/D vssd1 vssd1 vccd1 vccd1 _12367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11318_ vssd1 vssd1 vccd1 vccd1 _11318_/HI _11318_/LO sky130_fd_sc_hd__conb_1
X_12298_ _12558_/CLK _12298_/D vssd1 vssd1 vccd1 vccd1 _12298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11249_ vssd1 vssd1 vccd1 vccd1 _11249_/HI _11249_/LO sky130_fd_sc_hd__conb_1
XFILLER_45_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06790_ _06787_/X _06788_/X _12022_/X _06789_/X vssd1 vssd1 vccd1 vccd1 _06790_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08460_ _13052_/Q _10346_/B _13047_/Q _10331_/A _08459_/X vssd1 vssd1 vccd1 vccd1
+ _08474_/B sky130_fd_sc_hd__a221o_1
XFILLER_24_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07411_ _07474_/A vssd1 vssd1 vccd1 vccd1 _07459_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_17_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08391_ _08405_/A vssd1 vssd1 vccd1 vccd1 _08391_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_90_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07342_ _11442_/X _07338_/X _13066_/Q _07339_/X vssd1 vssd1 vccd1 vccd1 _13066_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07273_ _11551_/X _07263_/X _13086_/Q _07264_/X vssd1 vssd1 vccd1 vccd1 _13086_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09012_ _09016_/A _09016_/B _11642_/X vssd1 vssd1 vccd1 vccd1 _12586_/D sky130_fd_sc_hd__and3_1
X_06224_ _06044_/Y _06223_/Y _06044_/Y _06223_/Y vssd1 vssd1 vccd1 vccd1 _06224_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_191_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06155_ _12747_/Q _12715_/Q _06151_/Y _06154_/Y vssd1 vssd1 vccd1 vccd1 _06155_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_104_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06086_ _12728_/Q _12696_/Q _12728_/Q _12696_/Q vssd1 vssd1 vccd1 vccd1 _06091_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_105_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09914_ _12662_/Q vssd1 vssd1 vccd1 vccd1 _09914_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09845_ _06466_/Y _09844_/X _06466_/Y _09844_/X vssd1 vssd1 vccd1 vccd1 _09845_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_6_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09776_ _13219_/Q _13218_/Q _06603_/Y _06607_/Y vssd1 vssd1 vccd1 vccd1 _09777_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06988_ _11884_/X vssd1 vssd1 vccd1 vccd1 _06995_/A sky130_fd_sc_hd__inv_2
XFILLER_37_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08727_ _08729_/A vssd1 vssd1 vccd1 vccd1 _08727_/X sky130_fd_sc_hd__clkbuf_1
XPHY_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08658_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08669_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _07609_/A _07609_/B vssd1 vssd1 vccd1 vccd1 _12974_/D sky130_fd_sc_hd__nor2_1
XPHY_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08591_/A vssd1 vssd1 vccd1 vccd1 _08589_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10620_ _10620_/A vssd1 vssd1 vccd1 vccd1 _10620_/Y sky130_fd_sc_hd__inv_2
XPHY_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10551_ _11357_/X _10554_/B vssd1 vssd1 vccd1 vccd1 _10551_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13270_ _13286_/CLK _13270_/D _06267_/X vssd1 vssd1 vccd1 vccd1 _13270_/Q sky130_fd_sc_hd__dfrtp_1
X_10482_ _10482_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _10484_/B sky130_fd_sc_hd__nor2_2
XFILLER_194_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12221_ _06305_/X _13156_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12221_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ _10005_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12152_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11103_ _10742_/X _11071_/X _06368_/X _11058_/A _11072_/X vssd1 vssd1 vccd1 vccd1
+ _11103_/X sky130_fd_sc_hd__a221o_1
XFILLER_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12083_ _12082_/X _12447_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12083_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11034_ _11034_/A vssd1 vssd1 vccd1 vccd1 _11034_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12985_ _12985_/CLK _12985_/D vssd1 vssd1 vccd1 vccd1 _12985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11936_ _09586_/Y _12797_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11936_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11867_ _10175_/X _12810_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11867_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10818_ _12515_/Q _12327_/Q _12515_/Q _12327_/Q vssd1 vssd1 vccd1 vccd1 _10821_/B
+ sky130_fd_sc_hd__o2bb2ai_2
XPHY_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11798_ _11797_/X _12060_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12439_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10749_ _10736_/X _10746_/X _06365_/X _07008_/X _10747_/X vssd1 vssd1 vccd1 vccd1
+ _10749_/X sky130_fd_sc_hd__a221o_1
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12419_ _12430_/CLK _12419_/D vssd1 vssd1 vccd1 vccd1 _12419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07960_ _07800_/X _11485_/X _07962_/S vssd1 vssd1 vccd1 vccd1 _12896_/D sky130_fd_sc_hd__mux2_1
XFILLER_68_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06911_ _06899_/X _06903_/X _06904_/X vssd1 vssd1 vccd1 vccd1 _06911_/X sky130_fd_sc_hd__a21bo_1
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07891_ _10324_/A _11492_/S _07891_/C vssd1 vssd1 vccd1 vccd1 _07951_/A sky130_fd_sc_hd__or3_1
X_09630_ _09630_/A _09630_/B _09625_/A vssd1 vssd1 vccd1 vccd1 _09632_/B sky130_fd_sc_hd__or3b_4
XFILLER_68_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06842_ _06719_/X _06834_/X _06840_/Y _06841_/X _13193_/Q vssd1 vssd1 vccd1 vccd1
+ _13193_/D sky130_fd_sc_hd__a32o_1
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06773_ _12029_/X _06731_/X _12029_/X _06731_/X vssd1 vssd1 vccd1 vccd1 _06778_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09561_ _13180_/Q vssd1 vssd1 vccd1 vccd1 _09578_/A sky130_fd_sc_hd__inv_2
XFILLER_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08512_ _08504_/X _12254_/X _08499_/X _12764_/Q vssd1 vssd1 vccd1 vccd1 _12764_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09492_ _09492_/A vssd1 vssd1 vccd1 vccd1 _09492_/X sky130_fd_sc_hd__clkbuf_4
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08443_ _08441_/Y _10397_/A _08442_/Y _12895_/Q vssd1 vssd1 vccd1 vccd1 _08443_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ _08374_/A vssd1 vssd1 vccd1 vccd1 _08374_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07325_ _11449_/X _07321_/X _13073_/Q _07324_/X vssd1 vssd1 vccd1 vccd1 _13073_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07256_ _07266_/A vssd1 vssd1 vccd1 vccd1 _07256_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06207_ _13281_/Q vssd1 vssd1 vccd1 vccd1 _06207_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07187_ _11518_/X _07176_/X _13117_/Q _07177_/X vssd1 vssd1 vccd1 vccd1 _13117_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06138_ _12740_/Q _12708_/Q _06137_/X vssd1 vssd1 vccd1 vccd1 _06138_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06069_ _06069_/A _06068_/X vssd1 vssd1 vccd1 vccd1 _06182_/B sky130_fd_sc_hd__or2b_1
XFILLER_154_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09828_ _09804_/Y _09848_/A _09827_/Y vssd1 vssd1 vccd1 vccd1 _09828_/X sky130_fd_sc_hd__o21a_1
XFILLER_171_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09759_ _13216_/Q _09758_/A _06626_/Y _09758_/Y vssd1 vssd1 vccd1 vccd1 _09759_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _13241_/CLK _12770_/D _08496_/X vssd1 vssd1 vccd1 vccd1 _12770_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11721_ _10655_/X _11909_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12449_/D sky130_fd_sc_hd__mux2_1
XPHY_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11652_ _10537_/Y _10534_/Y _11704_/S vssd1 vssd1 vccd1 vccd1 _12364_/D sky130_fd_sc_hd__mux2_1
XPHY_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10603_ _10603_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _10603_/X sky130_fd_sc_hd__or2_1
XPHY_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11583_ _10417_/Y _09186_/A _11592_/S vssd1 vssd1 vccd1 vccd1 _11583_/X sky130_fd_sc_hd__mux2_1
XPHY_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10534_ _11361_/X vssd1 vssd1 vccd1 vccd1 _10534_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13253_ _13253_/CLK _13253_/D _06360_/X vssd1 vssd1 vccd1 vccd1 _13253_/Q sky130_fd_sc_hd__dfrtp_2
X_10465_ _08128_/X _10462_/Y _10459_/X _10467_/C vssd1 vssd1 vccd1 vccd1 _10465_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ _12203_/X _12622_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12204_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10396_ _10395_/A _10395_/B _10387_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10396_/Y
+ sky130_fd_sc_hd__a211oi_4
X_13184_ _13190_/CLK _13184_/D _06916_/X vssd1 vssd1 vccd1 vccd1 _13184_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ _12134_/X _12435_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12135_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12066_ _12445_/Q _10681_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _12066_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11017_ _12358_/Q _11018_/C _12358_/Q _11018_/C vssd1 vssd1 vccd1 vccd1 _12358_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ _12974_/CLK _12968_/D vssd1 vssd1 vccd1 vccd1 _12968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_66_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12973_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11919_ _11918_/X _12442_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _11919_/X sky130_fd_sc_hd__mux2_1
XPHY_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _12166_/X _12899_/D _07953_/X vssd1 vssd1 vccd1 vccd1 _12899_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07110_ _08271_/A _09978_/B _09296_/A vssd1 vssd1 vccd1 vccd1 _11522_/S sky130_fd_sc_hd__nor3_4
X_08090_ _08098_/A vssd1 vssd1 vccd1 vccd1 _08090_/X sky130_fd_sc_hd__clkbuf_1
X_07041_ _07059_/A vssd1 vssd1 vccd1 vccd1 _07042_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_173_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08992_ _12597_/Q vssd1 vssd1 vccd1 vccd1 _08992_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07943_ _07945_/A vssd1 vssd1 vccd1 vccd1 _07943_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07874_ _10368_/B vssd1 vssd1 vccd1 vccd1 _10362_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09613_ _13158_/Q _09475_/X _09598_/Y _09919_/B _09612_/X vssd1 vssd1 vccd1 vccd1
+ _09613_/Y sky130_fd_sc_hd__o221ai_2
X_06825_ _08854_/A vssd1 vssd1 vccd1 vccd1 _07477_/A sky130_fd_sc_hd__buf_4
XFILLER_44_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09544_ _12868_/Q vssd1 vssd1 vccd1 vccd1 _09544_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06756_ _11996_/X _06756_/B vssd1 vssd1 vccd1 vccd1 _06756_/X sky130_fd_sc_hd__or2_2
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06687_ _06690_/A vssd1 vssd1 vccd1 vccd1 _06687_/X sky130_fd_sc_hd__clkbuf_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09475_ _09475_/A vssd1 vssd1 vccd1 vccd1 _09475_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08426_ _12778_/Q _08417_/X _08005_/X _08418_/X vssd1 vssd1 vccd1 vccd1 _12778_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08357_ _08359_/A vssd1 vssd1 vccd1 vccd1 _08374_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07308_ _09185_/D vssd1 vssd1 vccd1 vccd1 _09226_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_109_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08288_ _12832_/Q _11607_/X _08292_/S vssd1 vssd1 vccd1 vccd1 _12832_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07239_ _07251_/A vssd1 vssd1 vccd1 vccd1 _07239_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_125_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10250_ _10248_/Y _10032_/X _10249_/Y _10028_/X vssd1 vssd1 vccd1 vccd1 _10250_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10181_ _12779_/Q vssd1 vssd1 vccd1 vccd1 _10181_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput580 _12297_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput591 _12563_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_121_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12822_ _12169_/X _12822_/D _08311_/X vssd1 vssd1 vccd1 vccd1 _12822_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12753_ _12753_/CLK _12753_/D _08543_/X vssd1 vssd1 vccd1 vccd1 _12753_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11703_/X _11889_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12394_/D sky130_fd_sc_hd__mux2_1
XPHY_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12685_/CLK _12684_/D _08744_/X vssd1 vssd1 vccd1 vccd1 _12684_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ _10505_/Y _12988_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11635_/X sky130_fd_sc_hd__mux2_1
XPHY_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ _12823_/Q _09180_/C _11569_/S vssd1 vssd1 vccd1 vccd1 _11566_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10517_ _12591_/Q _07765_/B _07766_/B vssd1 vssd1 vccd1 vccd1 _10517_/X sky130_fd_sc_hd__a21bo_1
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11497_ _10360_/Y _10528_/B _11501_/S vssd1 vssd1 vccd1 vccd1 _11497_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_113_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 _12707_/CLK sky130_fd_sc_hd__clkbuf_16
X_13236_ _13236_/CLK _13236_/D _06433_/X vssd1 vssd1 vccd1 vccd1 _13236_/Q sky130_fd_sc_hd__dfrtp_4
X_10448_ _10449_/B _10455_/D _12820_/Q _10447_/B _10437_/X vssd1 vssd1 vccd1 vccd1
+ _10448_/X sky130_fd_sc_hd__o221a_1
XFILLER_123_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13167_ _13170_/CLK _13167_/D _07022_/X vssd1 vssd1 vccd1 vccd1 _13167_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10379_ _10380_/B _10380_/C _12915_/Q _10377_/A _10350_/X vssd1 vssd1 vccd1 vccd1
+ _10379_/X sky130_fd_sc_hd__o221a_1
X_12118_ _12436_/Q _12117_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12118_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13098_ _12167_/X _13098_/D _07241_/X vssd1 vssd1 vccd1 vccd1 _13098_/Q sky130_fd_sc_hd__dfrtp_1
X_12049_ _10765_/Y _11122_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12049_/X sky130_fd_sc_hd__mux2_2
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06610_ _11894_/X _11892_/X _06609_/X vssd1 vssd1 vccd1 vccd1 _06610_/X sky130_fd_sc_hd__o21a_1
X_07590_ _07590_/A _12600_/Q vssd1 vssd1 vccd1 vccd1 _09276_/C sky130_fd_sc_hd__or2_4
XFILLER_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06541_ _12172_/X _11135_/A _06539_/X vssd1 vssd1 vccd1 vccd1 _06541_/X sky130_fd_sc_hd__a21bo_1
XFILLER_34_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09260_ _09029_/B _09288_/B _07508_/Y _08984_/Y vssd1 vssd1 vccd1 vccd1 _09260_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06472_ _11883_/X _10787_/A _11883_/X _10787_/A vssd1 vssd1 vccd1 vccd1 _06479_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08211_ _13084_/Q _08177_/Y _13107_/Q _08154_/Y vssd1 vssd1 vccd1 vccd1 _08211_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09191_ _09215_/A vssd1 vssd1 vccd1 vccd1 _09216_/A sky130_fd_sc_hd__inv_2
XFILLER_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08142_ _12805_/Q vssd1 vssd1 vccd1 vccd1 _10405_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08073_ _08085_/A vssd1 vssd1 vccd1 vccd1 _08073_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07024_ _07024_/A vssd1 vssd1 vccd1 vccd1 _07024_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput308 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _07097_/B sky130_fd_sc_hd__clkbuf_1
X_08975_ _09279_/C _12605_/Q _12600_/Q vssd1 vssd1 vccd1 vccd1 _08976_/B sky130_fd_sc_hd__a21oi_1
XFILLER_29_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput319 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 _07102_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07926_ _12910_/Q _11499_/X _07932_/S vssd1 vssd1 vccd1 vccd1 _12910_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07857_ _13023_/Q _10357_/B _13037_/Q _10393_/A vssd1 vssd1 vccd1 vccd1 _07857_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_57_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06808_ _11881_/X vssd1 vssd1 vccd1 vccd1 _06808_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07788_ _07566_/X _07780_/A _12927_/Q _07781_/A _07522_/A vssd1 vssd1 vccd1 vccd1
+ _12927_/D sky130_fd_sc_hd__a221o_1
XFILLER_45_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09527_ _09526_/A _09526_/B _09526_/C vssd1 vssd1 vccd1 vccd1 _09528_/B sky130_fd_sc_hd__o21a_1
X_06739_ _13204_/Q vssd1 vssd1 vccd1 vccd1 _06739_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _12982_/Q _09436_/A _12998_/Q _09451_/X vssd1 vssd1 vccd1 vccd1 _09458_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08409_ _12785_/Q _08401_/X _07983_/X _08403_/X vssd1 vssd1 vccd1 vccd1 _12785_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09389_ _12416_/D vssd1 vssd1 vccd1 vccd1 _10610_/B sky130_fd_sc_hd__inv_2
XFILLER_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11420_ _12895_/Q _09185_/C _11422_/S vssd1 vssd1 vccd1 vccd1 _11420_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11351_ _09453_/X _12988_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _12315_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10302_ _12652_/Q vssd1 vssd1 vccd1 vccd1 _10302_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11282_ vssd1 vssd1 vccd1 vccd1 _11282_/HI _11282_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13021_ _12164_/X _13021_/D _07463_/X vssd1 vssd1 vccd1 vccd1 _13021_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10233_ _12855_/Q vssd1 vssd1 vccd1 vccd1 _10233_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10164_ _12628_/Q vssd1 vssd1 vccd1 vccd1 _10164_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10095_ _12625_/Q vssd1 vssd1 vccd1 vccd1 _10095_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ _12169_/X _12805_/D _08350_/X vssd1 vssd1 vccd1 vccd1 _12805_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_188_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10997_ _10997_/A vssd1 vssd1 vccd1 vccd1 _10997_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12736_ _12737_/CLK _12736_/D _08613_/X vssd1 vssd1 vccd1 vccd1 _12736_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_71_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _12718_/CLK _12667_/D _08803_/X vssd1 vssd1 vccd1 vccd1 _12667_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ _12972_/Q _12985_/Q _12601_/Q vssd1 vssd1 vccd1 vccd1 _11618_/X sky130_fd_sc_hd__mux2_1
X_12598_ _12975_/CLK _12598_/D vssd1 vssd1 vccd1 vccd1 _12598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11549_ _12806_/Q _09185_/C _11550_/S vssd1 vssd1 vccd1 vccd1 _11549_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13219_ _13219_/CLK _13219_/D _06601_/X vssd1 vssd1 vccd1 vccd1 _13219_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12716_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08760_ _08781_/A vssd1 vssd1 vccd1 vccd1 _08760_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_81_wb_clk_i _12960_/CLK vssd1 vssd1 vccd1 vccd1 _13249_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07711_ _07711_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07711_/Y sky130_fd_sc_hd__nor2_1
X_08691_ _08699_/A vssd1 vssd1 vccd1 vccd1 _08691_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_10_wb_clk_i _12328_/CLK vssd1 vssd1 vccd1 vccd1 _12517_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07642_ _07665_/A _07642_/B _07666_/A vssd1 vssd1 vccd1 vccd1 _07654_/A sky130_fd_sc_hd__nor3_4
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07573_ _07575_/A vssd1 vssd1 vccd1 vccd1 _07574_/A sky130_fd_sc_hd__inv_2
XFILLER_20_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09312_ _09312_/A vssd1 vssd1 vccd1 vccd1 _12101_/S sky130_fd_sc_hd__inv_2
X_06524_ _06766_/A vssd1 vssd1 vccd1 vccd1 _06580_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09243_ _09243_/A _10528_/C _09243_/C _09243_/D vssd1 vssd1 vccd1 vccd1 _09245_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06455_ _06440_/X _06441_/Y _06420_/X _06454_/X vssd1 vssd1 vccd1 vccd1 _13235_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06386_ _13246_/Q vssd1 vssd1 vccd1 vccd1 _06386_/X sky130_fd_sc_hd__buf_2
X_09174_ _11619_/X _09163_/A _12494_/Q _09164_/A vssd1 vssd1 vccd1 vccd1 _12494_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08125_ _13120_/Q _10420_/A _08121_/Y _12814_/Q _08124_/X vssd1 vssd1 vccd1 vccd1
+ _08132_/C sky130_fd_sc_hd__a221o_1
XFILLER_179_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08056_ _12864_/Q _08040_/A _07300_/X _08041_/A vssd1 vssd1 vccd1 vccd1 _12864_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07007_ _07007_/A vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_190_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput105 la_data_in[44] vssd1 vssd1 vccd1 vccd1 input105/X sky130_fd_sc_hd__buf_1
Xinput116 la_data_in[54] vssd1 vssd1 vccd1 vccd1 input116/X sky130_fd_sc_hd__buf_1
XFILLER_131_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput127 la_data_in[64] vssd1 vssd1 vccd1 vccd1 input127/X sky130_fd_sc_hd__buf_1
X_08958_ _12142_/S _11909_/S vssd1 vssd1 vccd1 vccd1 _12619_/D sky130_fd_sc_hd__and2_1
XFILLER_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput138 la_data_in[74] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_hd__buf_1
XFILLER_9_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput149 la_data_in[84] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_hd__buf_1
XFILLER_76_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07909_ _07917_/A vssd1 vssd1 vccd1 vccd1 _07909_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08889_ _08883_/X _06295_/Y _08878_/X _12633_/Q vssd1 vssd1 vccd1 vccd1 _12633_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_186_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10920_ _10918_/Y _10919_/Y _12530_/Q _12342_/Q vssd1 vssd1 vccd1 vccd1 _10947_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_72_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10851_ _12520_/Q _12332_/Q _10849_/Y _10850_/Y vssd1 vssd1 vccd1 vccd1 _10851_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_147_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10782_/A vssd1 vssd1 vccd1 vccd1 _10782_/Y sky130_fd_sc_hd__inv_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12521_ _12802_/CLK _12521_/D vssd1 vssd1 vccd1 vccd1 _12521_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _12455_/CLK _12452_/D vssd1 vssd1 vccd1 vccd1 _12452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11403_ _10600_/X _12408_/D _11403_/S vssd1 vssd1 vccd1 vccd1 _11403_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12383_ _12472_/CLK _12383_/D vssd1 vssd1 vccd1 vccd1 _12405_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11334_ vssd1 vssd1 vccd1 vccd1 _11334_/HI _11334_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ vssd1 vssd1 vccd1 vccd1 _11265_/HI _11265_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13004_ _13004_/CLK _13004_/D vssd1 vssd1 vccd1 vccd1 _13004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10216_ _12854_/Q vssd1 vssd1 vccd1 vccd1 _10216_/Y sky130_fd_sc_hd__inv_2
X_11196_ vssd1 vssd1 vccd1 vccd1 _11196_/HI _11196_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _10142_/Y _10020_/X _10143_/Y _10018_/X _10146_/X vssd1 vssd1 vccd1 vccd1
+ _10147_/X sky130_fd_sc_hd__o221a_1
XFILLER_94_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10078_ _13149_/Q vssd1 vssd1 vccd1 vccd1 _10078_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12719_ _12719_/CLK _12719_/D _08653_/X vssd1 vssd1 vccd1 vccd1 _12719_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06240_ _13275_/Q vssd1 vssd1 vccd1 vccd1 _06240_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06171_ _06046_/A _06046_/B _06170_/X _06149_/Y vssd1 vssd1 vccd1 vccd1 _06171_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_144_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_1_wb_clk_i clkbuf_2_0_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09930_ _09928_/Y _09922_/X _06291_/A _09915_/X _09929_/X vssd1 vssd1 vccd1 vccd1
+ _09930_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_172_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09861_ _09492_/X _09859_/Y _09860_/X _09700_/A vssd1 vssd1 vccd1 vccd1 _09861_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_98_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08812_ _08798_/X _08801_/X _06300_/Y _12664_/Q _08811_/X vssd1 vssd1 vccd1 vccd1
+ _12664_/D sky130_fd_sc_hd__a32o_1
XFILLER_85_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09792_ _09792_/A vssd1 vssd1 vccd1 vccd1 _09802_/B sky130_fd_sc_hd__inv_2
XFILLER_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08743_ _08739_/Y _08565_/X _11963_/S _08742_/X vssd1 vssd1 vccd1 vccd1 _12685_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08674_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07625_ _12961_/Q _12960_/Q _12959_/Q _12958_/Q vssd1 vssd1 vccd1 vccd1 _07664_/A
+ sky130_fd_sc_hd__or4_4
XPHY_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07556_ _07775_/A vssd1 vssd1 vccd1 vccd1 _07556_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06507_ _06658_/A vssd1 vssd1 vccd1 vccd1 _06507_/X sky130_fd_sc_hd__buf_2
XFILLER_179_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07487_ _07489_/A vssd1 vssd1 vccd1 vccd1 _07487_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09226_ _09226_/A _09226_/B vssd1 vssd1 vccd1 vccd1 _09228_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06438_ _06465_/A vssd1 vssd1 vccd1 vccd1 _06438_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_166_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09157_ _11634_/X _09154_/X _12509_/Q _09156_/X vssd1 vssd1 vccd1 vccd1 _12509_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06369_ _06361_/X _12228_/X _06358_/X _06368_/X vssd1 vssd1 vccd1 vccd1 _13251_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_135_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08108_ _12834_/Q vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__clkbuf_2
X_09088_ _09123_/A vssd1 vssd1 vccd1 vccd1 _09115_/A sky130_fd_sc_hd__buf_4
XFILLER_123_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08039_ _08051_/A vssd1 vssd1 vccd1 vccd1 _08039_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11050_ _13241_/Q _11107_/A _10696_/A _06917_/A _06470_/Y vssd1 vssd1 vccd1 vccd1
+ _11099_/A sky130_fd_sc_hd__o221a_1
XFILLER_150_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10001_ _10001_/A vssd1 vssd1 vccd1 vccd1 _10001_/X sky130_fd_sc_hd__buf_2
XFILLER_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11952_ _09833_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11952_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _10903_/A vssd1 vssd1 vccd1 vccd1 _10921_/B sky130_fd_sc_hd__inv_2
XFILLER_199_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11883_ _10734_/X _10789_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _11883_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10834_ _12516_/Q _12328_/Q _10830_/X _12517_/Q _12329_/Q vssd1 vssd1 vccd1 vccd1
+ _10834_/X sky130_fd_sc_hd__a32o_1
XFILLER_198_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10765_ _10765_/A vssd1 vssd1 vccd1 vccd1 _10765_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ _13244_/CLK _12504_/D vssd1 vssd1 vccd1 vccd1 _12504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10696_ _10696_/A vssd1 vssd1 vccd1 vccd1 _10696_/X sky130_fd_sc_hd__buf_2
XFILLER_201_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12435_ _12441_/CLK _12435_/D vssd1 vssd1 vccd1 vccd1 _12435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12366_ _12369_/CLK _12366_/D vssd1 vssd1 vccd1 vccd1 _12366_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput409 _11191_/LO vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11317_ vssd1 vssd1 vccd1 vccd1 _11317_/HI _11317_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12297_ _12558_/CLK _12297_/D vssd1 vssd1 vccd1 vccd1 _12297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11248_ vssd1 vssd1 vccd1 vccd1 _11248_/HI _11248_/LO sky130_fd_sc_hd__conb_1
XFILLER_122_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ vssd1 vssd1 vccd1 vccd1 _11179_/HI _11179_/LO sky130_fd_sc_hd__conb_1
XFILLER_171_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07410_ _12843_/Q _11459_/S vssd1 vssd1 vccd1 vccd1 _07474_/A sky130_fd_sc_hd__or2_1
XFILLER_90_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08390_ _12791_/Q _08374_/A _07300_/X _08375_/A vssd1 vssd1 vccd1 vccd1 _12791_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07341_ _07345_/A vssd1 vssd1 vccd1 vccd1 _07341_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07272_ _07280_/A vssd1 vssd1 vccd1 vccd1 _07272_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09011_ _09016_/A _09016_/B _11643_/X vssd1 vssd1 vccd1 vccd1 _12587_/D sky130_fd_sc_hd__and3_1
X_06223_ _06041_/Y _06042_/Y _06145_/X _06045_/A vssd1 vssd1 vccd1 vccd1 _06223_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_191_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06154_ _06154_/A vssd1 vssd1 vccd1 vccd1 _06154_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06085_ _06180_/A _06180_/B vssd1 vssd1 vccd1 vccd1 _06132_/B sky130_fd_sc_hd__or2_1
XFILLER_105_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09913_ _12661_/Q _12611_/Q _06316_/X _09547_/A _09912_/Y vssd1 vssd1 vccd1 vccd1
+ _09913_/X sky130_fd_sc_hd__a221o_1
XFILLER_144_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09844_ _06483_/Y _06488_/Y _09836_/Y _09837_/Y vssd1 vssd1 vccd1 vccd1 _09844_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09775_ _06647_/Y _06651_/Y _06626_/Y _09758_/Y vssd1 vssd1 vccd1 vccd1 _09779_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_101_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06987_ _11879_/X vssd1 vssd1 vccd1 vccd1 _06987_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08726_ _11825_/X _08715_/X _12691_/Q _08716_/X vssd1 vssd1 vccd1 vccd1 _12691_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _08657_/A vssd1 vssd1 vccd1 vccd1 _08731_/A sky130_fd_sc_hd__buf_2
XPHY_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _12974_/Q _07610_/A _07607_/Y vssd1 vssd1 vccd1 vccd1 _07609_/B sky130_fd_sc_hd__o21a_1
XPHY_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _11954_/X _08575_/X _12745_/Q _08578_/X vssd1 vssd1 vccd1 vccd1 _12745_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07539_ _12999_/Q _07531_/X _09185_/B _07532_/X _07538_/X vssd1 vssd1 vccd1 vccd1
+ _12999_/D sky130_fd_sc_hd__o221a_1
XPHY_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10550_ _11357_/X vssd1 vssd1 vccd1 vccd1 _10550_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09209_ _12480_/Q _09207_/X _09244_/B _09208_/X vssd1 vssd1 vccd1 vccd1 _12480_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10481_ _12832_/Q _10478_/Y _10459_/X _10482_/B vssd1 vssd1 vccd1 vccd1 _10481_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12220_ _12219_/X _12630_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12220_/X sky130_fd_sc_hd__mux2_2
XFILLER_136_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12151_ _10004_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12151_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11102_ _06362_/X _11045_/A _08535_/A _10730_/X _07030_/X vssd1 vssd1 vccd1 vccd1
+ _11102_/X sky130_fd_sc_hd__a32o_1
X_12082_ _12447_/Q _12081_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _12082_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11033_ _11033_/A vssd1 vssd1 vccd1 vccd1 _11033_/X sky130_fd_sc_hd__buf_2
XFILLER_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_138_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _12870_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12984_ _12984_/CLK _12984_/D vssd1 vssd1 vccd1 vccd1 _12984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11935_ _09571_/X _12796_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11935_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11866_ _10150_/Y _12318_/Q _12312_/Q vssd1 vssd1 vccd1 vccd1 _11866_/X sky130_fd_sc_hd__mux2_2
XPHY_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10817_ _10821_/C _10821_/A _10821_/C _10821_/A vssd1 vssd1 vccd1 vccd1 _12326_/D
+ sky130_fd_sc_hd__a2bb2oi_1
XPHY_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11797_ _12060_/X _11796_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11797_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10748_ _10730_/X _10746_/X _06362_/X _07008_/X _10747_/X vssd1 vssd1 vccd1 vccd1
+ _10748_/X sky130_fd_sc_hd__a221o_1
XFILLER_159_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10679_ _10792_/B _11818_/S vssd1 vssd1 vccd1 vccd1 _10679_/X sky130_fd_sc_hd__and2_1
XFILLER_173_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12418_ _12430_/CLK _12418_/D vssd1 vssd1 vccd1 vccd1 _12418_/Q sky130_fd_sc_hd__dfxtp_1
X_12349_ _12537_/CLK _12349_/D vssd1 vssd1 vccd1 vccd1 _12349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06910_ _12003_/X _06896_/B _06896_/X vssd1 vssd1 vccd1 vccd1 _06910_/X sky130_fd_sc_hd__a21bo_1
XFILLER_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07890_ _07885_/Y _07887_/X _12840_/Q _07888_/Y _10054_/A vssd1 vssd1 vccd1 vccd1
+ _07891_/C sky130_fd_sc_hd__a221oi_2
XFILLER_110_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06841_ _06841_/A vssd1 vssd1 vccd1 vccd1 _06841_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09560_ _13154_/Q _09475_/X _09544_/Y _09919_/B _09559_/X vssd1 vssd1 vccd1 vccd1
+ _09560_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_110_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06772_ _06770_/X _06771_/X _06770_/X _06771_/X vssd1 vssd1 vccd1 vccd1 _06778_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08511_ _08518_/A vssd1 vssd1 vccd1 vccd1 _08511_/X sky130_fd_sc_hd__clkbuf_1
X_09491_ _09491_/A vssd1 vssd1 vccd1 vccd1 _09492_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08442_ _13044_/Q vssd1 vssd1 vccd1 vccd1 _08442_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ _08385_/A vssd1 vssd1 vccd1 vccd1 _08373_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07324_ _07369_/A vssd1 vssd1 vccd1 vccd1 _07324_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07255_ _11558_/X _07248_/X _13093_/Q _07249_/X vssd1 vssd1 vccd1 vccd1 _13093_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06206_ _06214_/A vssd1 vssd1 vccd1 vccd1 _06206_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07186_ _07206_/A vssd1 vssd1 vccd1 vccd1 _07186_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06137_ _12740_/Q _12708_/Q _12739_/Q _12707_/Q vssd1 vssd1 vccd1 vccd1 _06137_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06068_ _12734_/Q _12702_/Q _06067_/X vssd1 vssd1 vccd1 vccd1 _06068_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09827_ _09826_/Y _09800_/Y _09813_/X vssd1 vssd1 vccd1 vccd1 _09827_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09758_ _09758_/A vssd1 vssd1 vccd1 vccd1 _09758_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08709_ _11832_/X _08700_/X _12698_/Q _08701_/X vssd1 vssd1 vccd1 vccd1 _12698_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09689_ _13203_/Q vssd1 vssd1 vccd1 vccd1 _09689_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11719_/X _10652_/Y _11774_/S vssd1 vssd1 vccd1 vccd1 _12424_/D sky130_fd_sc_hd__mux2_1
XPHY_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _10532_/X _10532_/B _11704_/S vssd1 vssd1 vccd1 vccd1 _12363_/D sky130_fd_sc_hd__mux2_1
XPHY_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10602_ _10603_/B vssd1 vssd1 vccd1 vccd1 _10602_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11582_ _10414_/X _09186_/B _11610_/S vssd1 vssd1 vccd1 vccd1 _11582_/X sky130_fd_sc_hd__mux2_1
XPHY_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10533_ _12364_/Q _12363_/Q _09328_/B vssd1 vssd1 vccd1 vccd1 _10533_/Y sky130_fd_sc_hd__o21ai_1
XPHY_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13252_ _13252_/CLK _13252_/D _06364_/X vssd1 vssd1 vccd1 vccd1 _13252_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10464_ _10464_/A vssd1 vssd1 vccd1 vccd1 _10467_/C sky130_fd_sc_hd__inv_2
XFILLER_89_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12203_ _06351_/X _13147_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12203_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13183_ _13183_/CLK _13183_/D _06921_/X vssd1 vssd1 vccd1 vccd1 _13183_/Q sky130_fd_sc_hd__dfrtp_1
X_10395_ _10395_/A _10395_/B vssd1 vssd1 vccd1 vccd1 _10397_/B sky130_fd_sc_hd__nor2_4
XFILLER_159_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12134_ _12435_/Q _12133_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12134_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12065_ _12064_/X _12440_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12065_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11016_ _11018_/C _11016_/B vssd1 vssd1 vccd1 vccd1 _12357_/D sky130_fd_sc_hd__nor2_1
XFILLER_42_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12967_ _12974_/CLK _12967_/D vssd1 vssd1 vccd1 vccd1 _12967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11918_ _12442_/Q _11917_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _11918_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12898_ _12166_/X _12898_/D _07955_/X vssd1 vssd1 vccd1 vccd1 _12898_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11849_ _09960_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11849_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_35_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12415_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_147_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07040_ _07074_/A vssd1 vssd1 vccd1 vccd1 _07040_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08991_ _08988_/X _08990_/X _11147_/A vssd1 vssd1 vccd1 vccd1 _12600_/D sky130_fd_sc_hd__o21a_1
XFILLER_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07942_ _12903_/Q _11492_/X _07946_/S vssd1 vssd1 vccd1 vccd1 _12903_/D sky130_fd_sc_hd__mux2_1
XFILLER_141_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07873_ _12909_/Q vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__inv_2
X_09612_ _09952_/A _09949_/A _09611_/A _09611_/B _09623_/B vssd1 vssd1 vccd1 vccd1
+ _09612_/X sky130_fd_sc_hd__a221o_2
XFILLER_68_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06824_ _06824_/A vssd1 vssd1 vccd1 vccd1 _13196_/D sky130_fd_sc_hd__inv_2
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09543_ _09535_/Y _07069_/A _12867_/Q _07729_/X _09542_/X vssd1 vssd1 vccd1 vccd1
+ _09543_/X sky130_fd_sc_hd__a221o_1
X_06755_ _11993_/X vssd1 vssd1 vccd1 vccd1 _06756_/B sky130_fd_sc_hd__inv_2
XFILLER_3_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09474_ _09482_/A _09482_/B _13164_/Q _13163_/Q vssd1 vssd1 vccd1 vccd1 _09474_/X
+ sky130_fd_sc_hd__o22a_1
X_06686_ _06435_/X _12190_/X _06436_/X _13210_/Q vssd1 vssd1 vccd1 vccd1 _13210_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08425_ _08433_/A vssd1 vssd1 vccd1 vccd1 _08425_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _09969_/B _08399_/B vssd1 vssd1 vccd1 vccd1 _08359_/A sky130_fd_sc_hd__or2_1
XFILLER_165_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07307_ _07330_/A vssd1 vssd1 vccd1 vccd1 _07307_/X sky130_fd_sc_hd__clkbuf_1
X_08287_ _08296_/A vssd1 vssd1 vccd1 vccd1 _08287_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07238_ _07253_/A vssd1 vssd1 vccd1 vccd1 _07251_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07169_ _07477_/A vssd1 vssd1 vccd1 vccd1 _07253_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10180_ _10178_/Y _10000_/A _10179_/Y _10137_/X vssd1 vssd1 vccd1 vccd1 _10180_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput570 _11313_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput581 _12298_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput592 _12564_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12821_ _12169_/X _12821_/D _08314_/X vssd1 vssd1 vccd1 vccd1 _12821_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12752_ _12753_/CLK _12752_/D _08545_/X vssd1 vssd1 vccd1 vccd1 _12752_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11889_/X _09180_/A _11703_/S vssd1 vssd1 vccd1 vccd1 _11703_/X sky130_fd_sc_hd__mux2_1
XPHY_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12683_/CLK _12683_/D _08747_/X vssd1 vssd1 vccd1 vccd1 _12683_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_187_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _10504_/X _12933_/Q _11634_/S vssd1 vssd1 vccd1 vccd1 _11634_/X sky130_fd_sc_hd__mux2_1
XPHY_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11565_ _12822_/Q _09180_/D _11569_/S vssd1 vssd1 vccd1 vccd1 _11565_/X sky130_fd_sc_hd__mux2_1
XPHY_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10516_ _12590_/Q _07764_/B _07765_/B vssd1 vssd1 vccd1 vccd1 _10516_/X sky130_fd_sc_hd__a21bo_1
XFILLER_10_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11496_ _10356_/X _09243_/A _11501_/S vssd1 vssd1 vccd1 vccd1 _11496_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13235_ _13235_/CLK _13235_/D _06438_/X vssd1 vssd1 vccd1 vccd1 _13235_/Q sky130_fd_sc_hd__dfrtp_1
X_10447_ _10458_/A _10447_/B _10447_/C vssd1 vssd1 vccd1 vccd1 _10447_/Y sky130_fd_sc_hd__nor3_1
XFILLER_124_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13166_ _13170_/CLK _13166_/D _07024_/X vssd1 vssd1 vccd1 vccd1 _13166_/Q sky130_fd_sc_hd__dfrtp_1
X_10378_ _07815_/X _10375_/Y _10372_/X _10380_/C vssd1 vssd1 vccd1 vccd1 _10378_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12117_ _10674_/Y _12436_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12117_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_153_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12337_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13097_ _12167_/X _13097_/D _07243_/X vssd1 vssd1 vccd1 vccd1 _13097_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12048_ _10764_/X _11125_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12048_/X sky130_fd_sc_hd__mux2_2
XFILLER_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06540_ _12176_/X _12175_/X _06539_/X vssd1 vssd1 vccd1 vccd1 _06540_/X sky130_fd_sc_hd__o21a_1
X_06471_ _06356_/X _11107_/A _06427_/X _06917_/A _06470_/Y vssd1 vssd1 vccd1 vccd1
+ _10787_/A sky130_fd_sc_hd__o221a_2
XFILLER_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08210_ _13090_/Q vssd1 vssd1 vccd1 vccd1 _08210_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09190_ _09215_/A vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08141_ _13115_/Q vssd1 vssd1 vccd1 vccd1 _08141_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08072_ _08284_/A vssd1 vssd1 vccd1 vccd1 _08085_/A sky130_fd_sc_hd__buf_2
XFILLER_119_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07023_ _06663_/X _12184_/X _06415_/B _13167_/Q vssd1 vssd1 vccd1 vccd1 _13167_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_114_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08974_ _09008_/A _13000_/Q _12571_/Q vssd1 vssd1 vccd1 vccd1 _12606_/D sky130_fd_sc_hd__and3_1
Xinput309 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _07097_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07925_ _07931_/A vssd1 vssd1 vccd1 vccd1 _07925_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07856_ _13028_/Q _10367_/A _07855_/Y _12911_/Q vssd1 vssd1 vccd1 vccd1 _07858_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06807_ _11880_/X vssd1 vssd1 vccd1 vccd1 _06807_/Y sky130_fd_sc_hd__inv_2
X_07787_ _07564_/X _07780_/X _12928_/Q _07781_/X _07522_/A vssd1 vssd1 vccd1 vccd1
+ _12928_/D sky130_fd_sc_hd__a221o_1
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09526_ _09526_/A _09526_/B _09526_/C vssd1 vssd1 vccd1 vccd1 _09528_/A sky130_fd_sc_hd__nor3_4
X_06738_ _06750_/A vssd1 vssd1 vccd1 vccd1 _06738_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _12930_/Q _09438_/X _12970_/Q _09440_/X vssd1 vssd1 vccd1 vccd1 _09457_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_196_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06669_ _06666_/X _06667_/X _12052_/X _06668_/X vssd1 vssd1 vccd1 vccd1 _06669_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08408_ _08420_/A vssd1 vssd1 vccd1 vccd1 _08408_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09388_ _12399_/D vssd1 vssd1 vccd1 vccd1 _10520_/C sky130_fd_sc_hd__inv_2
XFILLER_200_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08339_ _08339_/A vssd1 vssd1 vccd1 vccd1 _08339_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11350_ _09449_/X _12987_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _12314_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10301_ _13161_/Q vssd1 vssd1 vccd1 vccd1 _10301_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11281_ vssd1 vssd1 vccd1 vccd1 _11281_/HI _11281_/LO sky130_fd_sc_hd__conb_1
XFILLER_152_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13020_ _12164_/X _13020_/D _07465_/X vssd1 vssd1 vccd1 vccd1 _13020_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10232_ _13265_/Q vssd1 vssd1 vccd1 vccd1 _10232_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10163_ _10163_/A vssd1 vssd1 vccd1 vccd1 _10163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10094_ _07795_/Y _10070_/X _10093_/X vssd1 vssd1 vccd1 vccd1 _10094_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12804_ _12169_/X _12804_/D _08352_/X vssd1 vssd1 vccd1 vccd1 _12804_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_16_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10996_ _12540_/Q _12352_/Q _10988_/Y _10991_/X vssd1 vssd1 vccd1 vccd1 _10997_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12735_ _12735_/CLK _12735_/D _08615_/X vssd1 vssd1 vccd1 vccd1 _12735_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_76_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _13268_/CLK _12666_/D _08805_/X vssd1 vssd1 vccd1 vccd1 _12666_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11617_ _12971_/Q _12984_/Q _12601_/Q vssd1 vssd1 vccd1 vccd1 _11617_/X sky130_fd_sc_hd__mux2_1
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _12975_/CLK _12597_/D vssd1 vssd1 vccd1 vccd1 _12597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11548_ _12805_/Q _09185_/D _11578_/S vssd1 vssd1 vccd1 vccd1 _11548_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11479_ _12922_/Q _10794_/A _11481_/S vssd1 vssd1 vccd1 vccd1 _11479_/X sky130_fd_sc_hd__mux2_1
X_13218_ _13223_/CLK _13218_/D _06606_/X vssd1 vssd1 vccd1 vccd1 _13218_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13149_ _13152_/CLK _13149_/D _07076_/X vssd1 vssd1 vccd1 vccd1 _13149_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_151_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07710_ _12308_/Q vssd1 vssd1 vccd1 vccd1 _07711_/A sky130_fd_sc_hd__inv_2
XFILLER_111_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08690_ _11840_/X _08685_/X _12706_/Q _08686_/X vssd1 vssd1 vccd1 vccd1 _12706_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07641_ _12957_/Q _07646_/D vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__or2_2
XFILLER_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07572_ _07778_/A _09439_/A vssd1 vssd1 vccd1 vccd1 _07575_/A sky130_fd_sc_hd__or2_2
XFILLER_80_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12995_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09311_ _09311_/A vssd1 vssd1 vccd1 vccd1 _12141_/S sky130_fd_sc_hd__inv_8
XFILLER_20_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06523_ _06435_/X _12192_/X _06436_/X _13226_/Q vssd1 vssd1 vccd1 vccd1 _13226_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09242_ _09242_/A vssd1 vssd1 vccd1 vccd1 _10528_/A sky130_fd_sc_hd__inv_2
X_06454_ _06444_/Y _06451_/A _06453_/Y vssd1 vssd1 vccd1 vccd1 _06454_/X sky130_fd_sc_hd__o21a_1
XFILLER_179_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09173_ _11620_/X _09163_/A _12495_/Q _09164_/A vssd1 vssd1 vccd1 vccd1 _12495_/D
+ sky130_fd_sc_hd__a22o_1
X_06385_ _06391_/A vssd1 vssd1 vccd1 vccd1 _06385_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08124_ _13145_/Q _08122_/Y _13127_/Q _10439_/A vssd1 vssd1 vccd1 vccd1 _08124_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08055_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08055_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_179_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07006_ _07006_/A vssd1 vssd1 vccd1 vccd1 _07006_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput106 la_data_in[45] vssd1 vssd1 vccd1 vccd1 input106/X sky130_fd_sc_hd__buf_1
XFILLER_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput117 la_data_in[55] vssd1 vssd1 vccd1 vccd1 input117/X sky130_fd_sc_hd__buf_1
XFILLER_102_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput128 la_data_in[65] vssd1 vssd1 vccd1 vccd1 input128/X sky130_fd_sc_hd__buf_1
X_08957_ _09304_/A _12449_/Q vssd1 vssd1 vccd1 vccd1 _11909_/S sky130_fd_sc_hd__nor2_8
Xinput139 la_data_in[75] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_hd__buf_1
XFILLER_130_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07908_ _12918_/Q _11507_/X _07918_/S vssd1 vssd1 vccd1 vccd1 _12918_/D sky130_fd_sc_hd__mux2_1
X_08888_ _08897_/A vssd1 vssd1 vccd1 vccd1 _08888_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07839_ _10352_/B vssd1 vssd1 vccd1 vccd1 _07839_/X sky130_fd_sc_hd__buf_1
XFILLER_186_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10850_ _12332_/Q vssd1 vssd1 vccd1 vccd1 _10850_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _09505_/Y _09506_/Y _09508_/X vssd1 vssd1 vccd1 vccd1 _09509_/Y sky130_fd_sc_hd__o21ai_1
X_10781_ _10781_/A vssd1 vssd1 vccd1 vccd1 _10781_/Y sky130_fd_sc_hd__inv_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12520_ _12550_/CLK _12520_/D vssd1 vssd1 vccd1 vccd1 _12520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12467_/CLK _12451_/D vssd1 vssd1 vccd1 vccd1 _12451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11402_ _10618_/X _12412_/D _11889_/S vssd1 vssd1 vccd1 vccd1 _11402_/X sky130_fd_sc_hd__mux2_1
X_12382_ _12410_/CLK _12382_/D vssd1 vssd1 vccd1 vccd1 _12404_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_197_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11333_ vssd1 vssd1 vccd1 vccd1 _11333_/HI _11333_/LO sky130_fd_sc_hd__conb_1
XFILLER_158_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11264_ vssd1 vssd1 vccd1 vccd1 _11264_/HI _11264_/LO sky130_fd_sc_hd__conb_1
XFILLER_106_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13003_ _13004_/CLK _13003_/D vssd1 vssd1 vccd1 vccd1 _13003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10215_ _13264_/Q vssd1 vssd1 vccd1 vccd1 _10215_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_11195_ vssd1 vssd1 vccd1 vccd1 _11195_/HI _11195_/LO sky130_fd_sc_hd__conb_1
XFILLER_121_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10146_ _10144_/Y _10023_/X _10145_/Y _10025_/X vssd1 vssd1 vccd1 vccd1 _10146_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10077_ _10075_/Y _10018_/X _10076_/Y _10020_/X vssd1 vssd1 vccd1 vccd1 _10088_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_130_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10979_ _10969_/Y _10970_/Y _10966_/Y _10977_/C _10978_/X vssd1 vssd1 vccd1 vccd1
+ _10980_/B sky130_fd_sc_hd__o221a_1
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12718_ _12718_/CLK _12718_/D _08659_/X vssd1 vssd1 vccd1 vccd1 _12718_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ _12653_/CLK _12649_/D _08846_/X vssd1 vssd1 vccd1 vccd1 _12649_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06170_ _06138_/Y _06209_/B _06147_/Y vssd1 vssd1 vccd1 vccd1 _06170_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09860_ _09860_/A _09866_/B vssd1 vssd1 vccd1 vccd1 _09860_/X sky130_fd_sc_hd__or2_1
XFILLER_124_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08811_ _08811_/A vssd1 vssd1 vccd1 vccd1 _08811_/X sky130_fd_sc_hd__clkbuf_2
X_09791_ _09780_/A _09790_/A _09780_/Y _09790_/Y vssd1 vssd1 vccd1 vccd1 _09792_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08742_ _08764_/A vssd1 vssd1 vccd1 vccd1 _08742_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08673_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08684_/A sky130_fd_sc_hd__clkbuf_2
XPHY_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07624_ _12952_/Q _12949_/Q vssd1 vssd1 vccd1 vccd1 _07658_/A sky130_fd_sc_hd__or2_4
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07555_ _07545_/X _07552_/X _12993_/Q _07553_/X _09002_/A vssd1 vssd1 vccd1 vccd1
+ _12993_/D sky130_fd_sc_hd__a221o_1
XPHY_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06506_ _06522_/A vssd1 vssd1 vccd1 vccd1 _06506_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07486_ _11453_/X _07474_/X _13012_/Q _07475_/X vssd1 vssd1 vccd1 vccd1 _13012_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09225_ _12467_/Q _09083_/A _10792_/B _09247_/A vssd1 vssd1 vccd1 vccd1 _12467_/D
+ sky130_fd_sc_hd__a22o_1
X_06437_ _06435_/X _12193_/X _06436_/X _13236_/Q vssd1 vssd1 vccd1 vccd1 _13236_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09156_ _09164_/A vssd1 vssd1 vccd1 vccd1 _09156_/X sky130_fd_sc_hd__clkbuf_2
X_06368_ _13251_/Q vssd1 vssd1 vccd1 vccd1 _06368_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08107_ _13144_/Q vssd1 vssd1 vccd1 vccd1 _08107_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09087_ _09087_/A _10527_/D vssd1 vssd1 vccd1 vccd1 _09123_/A sky130_fd_sc_hd__or2_2
X_06299_ _06091_/A _06298_/X _06091_/A _06298_/X vssd1 vssd1 vccd1 vccd1 _06300_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08038_ _08038_/A vssd1 vssd1 vccd1 vccd1 _08051_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10000_ _10000_/A vssd1 vssd1 vccd1 vccd1 _10000_/X sky130_fd_sc_hd__buf_2
XFILLER_7_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09989_ _09973_/Y _10141_/A _09979_/X _09988_/X vssd1 vssd1 vccd1 vccd1 _10001_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11951_ _09819_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11951_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10902_ _12526_/Q _12338_/Q _10895_/Y _10896_/Y vssd1 vssd1 vccd1 vccd1 _10904_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11882_ _11043_/X _11039_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _11882_/X sky130_fd_sc_hd__mux2_2
XFILLER_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10833_ _10831_/Y _10832_/Y _10831_/Y _10832_/Y vssd1 vssd1 vccd1 vccd1 _12329_/D
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10764_ _10763_/X _10759_/X _06379_/X _10760_/X _10761_/X vssd1 vssd1 vccd1 vccd1
+ _10764_/X sky130_fd_sc_hd__a221o_1
XFILLER_41_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12503_ _13244_/CLK _12503_/D vssd1 vssd1 vccd1 vccd1 _12503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10695_ _13241_/Q vssd1 vssd1 vccd1 vccd1 _10696_/A sky130_fd_sc_hd__inv_2
XFILLER_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12434_ _12434_/CLK _12434_/D vssd1 vssd1 vccd1 vccd1 _12434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12365_ _12422_/CLK _12365_/D vssd1 vssd1 vccd1 vccd1 _12365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11316_ vssd1 vssd1 vccd1 vccd1 _11316_/HI _11316_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12296_ _12296_/CLK _12296_/D vssd1 vssd1 vccd1 vccd1 _12296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11247_ vssd1 vssd1 vccd1 vccd1 _11247_/HI _11247_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11178_ vssd1 vssd1 vccd1 vccd1 _11178_/HI _11178_/LO sky130_fd_sc_hd__conb_1
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10129_ _10150_/A _11976_/X vssd1 vssd1 vccd1 vccd1 _10129_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07340_ _11443_/X _07338_/X _13067_/Q _07339_/X vssd1 vssd1 vccd1 vccd1 _13067_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07271_ _11552_/X _07263_/X _13087_/Q _07264_/X vssd1 vssd1 vccd1 vccd1 _13087_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09010_ _13001_/Q vssd1 vssd1 vccd1 vccd1 _09016_/B sky130_fd_sc_hd__buf_1
X_06222_ _13279_/Q vssd1 vssd1 vccd1 vccd1 _06222_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06153_ _12746_/Q _12714_/Q _06152_/X vssd1 vssd1 vccd1 vccd1 _06154_/A sky130_fd_sc_hd__o21ai_2
XFILLER_176_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06084_ _12729_/Q _12697_/Q _06082_/Y _06083_/Y vssd1 vssd1 vccd1 vccd1 _06180_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09912_ _12884_/Q _09919_/B vssd1 vssd1 vccd1 vccd1 _09912_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09843_ _09701_/X _09841_/Y _09842_/X _09700_/A vssd1 vssd1 vccd1 vccd1 _09843_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06986_ _13175_/Q vssd1 vssd1 vccd1 vccd1 _09552_/B sky130_fd_sc_hd__inv_2
X_09774_ _09756_/X _09759_/X _09755_/Y _09760_/X vssd1 vssd1 vccd1 vccd1 _09782_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08725_ _08729_/A vssd1 vssd1 vccd1 vccd1 _08725_/X sky130_fd_sc_hd__clkbuf_1
XPHY_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _11928_/X _08654_/X _12719_/Q _08655_/X vssd1 vssd1 vccd1 vccd1 _12719_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _12601_/Q _07598_/C _12974_/Q vssd1 vssd1 vccd1 vccd1 _07607_/Y sky130_fd_sc_hd__o21ai_1
XPHY_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _08591_/A vssd1 vssd1 vccd1 vccd1 _08587_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ _08978_/A vssd1 vssd1 vccd1 vccd1 _07538_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07469_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07469_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09208_ _09216_/A vssd1 vssd1 vccd1 vccd1 _09208_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10480_ _10480_/A _10480_/B vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__or2_2
XFILLER_183_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09139_ _12500_/Q _09139_/B vssd1 vssd1 vccd1 vccd1 _09140_/B sky130_fd_sc_hd__or2_1
XFILLER_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12150_ _10002_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12150_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11101_ _10699_/X _11100_/X _13242_/Q _10769_/X _10770_/X vssd1 vssd1 vccd1 vccd1
+ _11101_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12081_ _12447_/Q _12080_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _12081_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11032_ _12755_/Q vssd1 vssd1 vccd1 vccd1 _11032_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12983_ _12984_/CLK _12983_/D vssd1 vssd1 vccd1 vccd1 _12983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11934_ _09560_/Y _12795_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11934_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11865_ _10153_/Y _12809_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11865_/X sky130_fd_sc_hd__mux2_1
XPHY_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_107_wb_clk_i _12726_/CLK vssd1 vssd1 vccd1 vccd1 _12695_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10816_ _10814_/Y _10815_/Y _12514_/Q _12326_/Q vssd1 vssd1 vccd1 vccd1 _10821_/A
+ sky130_fd_sc_hd__a22o_2
X_11796_ _09243_/A _11795_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11796_/X sky130_fd_sc_hd__mux2_1
XPHY_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10747_ _11899_/X vssd1 vssd1 vccd1 vccd1 _10747_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10678_ _12439_/Q _09315_/A _12440_/Q vssd1 vssd1 vccd1 vccd1 _10678_/X sky130_fd_sc_hd__o21a_1
XFILLER_185_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12417_ _12430_/CLK _12417_/D vssd1 vssd1 vccd1 vccd1 _12417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ _12540_/CLK _12348_/D vssd1 vssd1 vccd1 vccd1 _12348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12279_ _10279_/X _12905_/Q _11875_/X _10275_/Y _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12295_/D sky130_fd_sc_hd__mux4_2
XFILLER_141_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06840_ _12031_/X _06840_/B vssd1 vssd1 vccd1 vccd1 _06840_/Y sky130_fd_sc_hd__nand2_2
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06771_ _06754_/A _06754_/B _06754_/X vssd1 vssd1 vccd1 vccd1 _06771_/X sky130_fd_sc_hd__a21bo_1
XFILLER_83_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08510_ _08504_/X _12256_/X _08499_/X _12765_/Q vssd1 vssd1 vccd1 vccd1 _12765_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09490_ _09490_/A _09490_/B vssd1 vssd1 vccd1 vccd1 _09504_/A sky130_fd_sc_hd__and2_1
XFILLER_64_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08441_ _13072_/Q vssd1 vssd1 vccd1 vccd1 _08441_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08372_ _08372_/A vssd1 vssd1 vccd1 vccd1 _08385_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07323_ _07385_/A vssd1 vssd1 vccd1 vccd1 _07369_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_182_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07254_ _07266_/A vssd1 vssd1 vccd1 vccd1 _07254_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06205_ _06203_/Y _06022_/X _06163_/X _06204_/X vssd1 vssd1 vccd1 vccd1 _13282_/D
+ sky130_fd_sc_hd__o22ai_1
X_07185_ _07253_/A vssd1 vssd1 vccd1 vccd1 _07206_/A sky130_fd_sc_hd__buf_2
XFILLER_118_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06136_ _12738_/Q _12706_/Q _06135_/X vssd1 vssd1 vccd1 vccd1 _06136_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_105_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06067_ _06067_/A _06067_/B vssd1 vssd1 vccd1 vccd1 _06067_/X sky130_fd_sc_hd__or2_1
XFILLER_132_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09826_ _09826_/A vssd1 vssd1 vccd1 vccd1 _09826_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09757_ _13215_/Q _13214_/Q _06647_/Y _06651_/Y vssd1 vssd1 vccd1 vccd1 _09758_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_5_wb_clk_i _12844_/CLK vssd1 vssd1 vccd1 vccd1 _13146_/CLK sky130_fd_sc_hd__clkbuf_16
X_06969_ _12054_/X _06945_/X _12054_/X _06945_/X vssd1 vssd1 vccd1 vccd1 _06977_/B
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_104_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08708_ _08714_/A vssd1 vssd1 vccd1 vccd1 _08708_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09688_ _13202_/Q _13201_/Q _06763_/Y _06768_/Y vssd1 vssd1 vccd1 vccd1 _09690_/A
+ sky130_fd_sc_hd__o22a_1
XPHY_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08685_/A vssd1 vssd1 vccd1 vccd1 _08639_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11649_/X _10526_/Y _11704_/S vssd1 vssd1 vccd1 vccd1 _12371_/D sky130_fd_sc_hd__mux2_1
XPHY_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10601_ _10607_/A _11403_/X vssd1 vssd1 vccd1 vccd1 _10601_/Y sky130_fd_sc_hd__nor2b_1
XPHY_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11581_ _10412_/Y _09185_/C _11610_/S vssd1 vssd1 vccd1 vccd1 _11581_/X sky130_fd_sc_hd__mux2_1
XPHY_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10532_ _10535_/A _10532_/B vssd1 vssd1 vccd1 vccd1 _10532_/X sky130_fd_sc_hd__and2_1
XPHY_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13251_ _13252_/CLK _13251_/D _06367_/X vssd1 vssd1 vccd1 vccd1 _13251_/Q sky130_fd_sc_hd__dfrtp_2
X_10463_ _12825_/Q _12824_/Q _10463_/C vssd1 vssd1 vccd1 vccd1 _10464_/A sky130_fd_sc_hd__and3_1
XFILLER_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12202_ _11133_/X _10777_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _12202_/X sky130_fd_sc_hd__mux2_2
XFILLER_170_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13182_ _13190_/CLK _13182_/D _06937_/X vssd1 vssd1 vccd1 vccd1 _13182_/Q sky130_fd_sc_hd__dfrtp_1
X_10394_ _12921_/Q _10391_/Y _10372_/X _10395_/B vssd1 vssd1 vccd1 vccd1 _10394_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12133_ _10673_/X _12435_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12133_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12064_ _12063_/X _12440_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12064_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11015_ _11013_/A _11010_/A _11013_/B vssd1 vssd1 vccd1 vccd1 _11016_/B sky130_fd_sc_hd__o21a_1
XFILLER_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12966_ _12973_/CLK _12966_/D vssd1 vssd1 vccd1 vccd1 _12966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11917_ _12442_/Q _11916_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _11917_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12166_/X _12897_/D _07957_/X vssd1 vssd1 vccd1 vccd1 _12897_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_61_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _09959_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11848_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11779_ _12136_/X _12479_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11779_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_75_wb_clk_i _13219_/CLK vssd1 vssd1 vccd1 vccd1 _13208_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08990_ _07661_/A _07689_/B _08989_/Y _12597_/Q vssd1 vssd1 vccd1 vccd1 _08990_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07941_ _07945_/A vssd1 vssd1 vccd1 vccd1 _07941_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07872_ _13038_/Q _10395_/A _13033_/Q _07868_/Y vssd1 vssd1 vccd1 vccd1 _07879_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_09611_ _09611_/A _09611_/B vssd1 vssd1 vccd1 vccd1 _09623_/B sky130_fd_sc_hd__nor2_1
X_06823_ _06658_/A _06813_/X _06821_/X _06646_/X _06822_/Y vssd1 vssd1 vccd1 vccd1
+ _06824_/A sky130_fd_sc_hd__a32o_1
XFILLER_55_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06754_ _06754_/A _06754_/B vssd1 vssd1 vccd1 vccd1 _06754_/X sky130_fd_sc_hd__or2_1
XFILLER_3_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09542_ _09528_/A _09530_/X _09540_/Y _09491_/A _09541_/Y vssd1 vssd1 vccd1 vccd1
+ _09542_/X sky130_fd_sc_hd__o311a_1
XFILLER_58_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06685_ _06690_/A vssd1 vssd1 vccd1 vccd1 _06685_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09473_ _13163_/Q vssd1 vssd1 vccd1 vccd1 _09482_/B sky130_fd_sc_hd__inv_2
XFILLER_93_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08424_ _12779_/Q _08417_/X _07545_/X _08418_/X vssd1 vssd1 vccd1 vccd1 _12779_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_196_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ _08370_/A vssd1 vssd1 vccd1 vccd1 _08355_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07306_ _07362_/A vssd1 vssd1 vccd1 vccd1 _07330_/A sky130_fd_sc_hd__buf_2
XFILLER_192_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08286_ _12833_/Q _11608_/X _08292_/S vssd1 vssd1 vccd1 vccd1 _12833_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07237_ _11565_/X _07233_/X _13100_/Q _07234_/X vssd1 vssd1 vccd1 vccd1 _13100_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07168_ _11525_/X _07160_/X _13124_/Q _07161_/X vssd1 vssd1 vccd1 vccd1 _13124_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06119_ _06117_/Y _06118_/Y _12719_/Q _12687_/Q vssd1 vssd1 vccd1 vccd1 _06122_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_106_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07099_ _09071_/A _09071_/B _07099_/C _09041_/B vssd1 vssd1 vccd1 vccd1 _07317_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput560 _11304_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput571 _11314_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput582 _12555_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput593 _12565_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09809_ _09701_/X _09807_/Y _09808_/X _09682_/X vssd1 vssd1 vccd1 vccd1 _09809_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12820_ _12169_/X _12820_/D _08316_/X vssd1 vssd1 vccd1 vccd1 _12820_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12751_ _12751_/CLK _12751_/D _08549_/X vssd1 vssd1 vccd1 vccd1 _12751_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11701_/X _11887_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12393_/D sky130_fd_sc_hd__mux2_1
XPHY_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12682_/CLK _12682_/D _08752_/X vssd1 vssd1 vccd1 vccd1 _12682_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _10503_/X _12932_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11633_/X sky130_fd_sc_hd__mux2_1
XPHY_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11564_ _12821_/Q _09179_/A _11569_/S vssd1 vssd1 vccd1 vccd1 _11564_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10515_ _12589_/Q _07763_/B _07764_/B vssd1 vssd1 vccd1 vccd1 _10515_/X sky130_fd_sc_hd__a21bo_1
XFILLER_144_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11495_ _10355_/Y input333/X _11501_/S vssd1 vssd1 vccd1 vccd1 _11495_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13234_ _13237_/CLK _13234_/D _06456_/X vssd1 vssd1 vccd1 vccd1 _13234_/Q sky130_fd_sc_hd__dfrtp_2
X_10446_ _10444_/B _10444_/C _10444_/A vssd1 vssd1 vccd1 vccd1 _10447_/C sky130_fd_sc_hd__o21a_1
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10377_ _10377_/A vssd1 vssd1 vccd1 vccd1 _10380_/C sky130_fd_sc_hd__inv_2
X_13165_ _13170_/CLK _13165_/D _07027_/X vssd1 vssd1 vccd1 vccd1 _13165_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12116_ _10710_/Y _06446_/B _12768_/Q vssd1 vssd1 vccd1 vccd1 _12116_/X sky130_fd_sc_hd__mux2_2
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13096_ _12167_/X _13096_/D _07245_/X vssd1 vssd1 vccd1 vccd1 _13096_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12047_ _10756_/X _11124_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _12047_/X sky130_fd_sc_hd__mux2_2
XFILLER_172_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_122_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 _12679_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12949_ _12955_/CLK _12949_/D vssd1 vssd1 vccd1 vccd1 _12949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06470_ _12132_/X vssd1 vssd1 vccd1 vccd1 _06470_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08140_ _13124_/Q _10433_/B _13119_/Q _10418_/A _08139_/X vssd1 vssd1 vccd1 vccd1
+ _08163_/B sky130_fd_sc_hd__a221o_1
XFILLER_144_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08071_ _12859_/Q _08066_/X _07980_/X _08068_/X vssd1 vssd1 vccd1 vccd1 _12859_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07022_ _07024_/A vssd1 vssd1 vccd1 vccd1 _07022_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08973_ _09009_/A vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07924_ _12911_/Q _11500_/X _07932_/S vssd1 vssd1 vccd1 vccd1 _12911_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07855_ _13027_/Q vssd1 vssd1 vccd1 vccd1 _07855_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06806_ _06806_/A vssd1 vssd1 vccd1 vccd1 _06806_/X sky130_fd_sc_hd__clkbuf_1
X_07786_ _07562_/X _07780_/X _12929_/Q _07781_/X _07775_/X vssd1 vssd1 vccd1 vccd1
+ _12929_/D sky130_fd_sc_hd__a221o_1
X_09525_ _09524_/A _09524_/B _09524_/Y vssd1 vssd1 vccd1 vccd1 _09526_/C sky130_fd_sc_hd__a21o_1
X_06737_ _06737_/A vssd1 vssd1 vccd1 vccd1 _13205_/D sky130_fd_sc_hd__inv_2
XFILLER_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_52_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06668_ _06666_/X _06667_/X _06666_/X _06667_/X vssd1 vssd1 vccd1 vccd1 _06668_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09456_ _12969_/Q _09440_/X _09454_/X _09455_/X vssd1 vssd1 vccd1 vccd1 _09456_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08407_ _08521_/A vssd1 vssd1 vccd1 vccd1 _08420_/A sky130_fd_sc_hd__buf_2
XFILLER_101_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09387_ _12455_/Q _10599_/A _09366_/Y _12399_/D _09386_/X vssd1 vssd1 vccd1 vccd1
+ _09402_/A sky130_fd_sc_hd__o221a_1
XFILLER_71_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06599_ _06507_/X _06581_/Y _06489_/X _06598_/Y vssd1 vssd1 vccd1 vccd1 _13220_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08338_ _08117_/X _11586_/X _08349_/S vssd1 vssd1 vccd1 vccd1 _12811_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08269_ _13080_/Q vssd1 vssd1 vccd1 vccd1 _08269_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ _12636_/Q vssd1 vssd1 vccd1 vccd1 _10300_/Y sky130_fd_sc_hd__inv_2
X_11280_ vssd1 vssd1 vccd1 vccd1 _11280_/HI _11280_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10231_ _13018_/Q _10228_/X _13051_/Q _10229_/X vssd1 vssd1 vccd1 vccd1 _10231_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10162_ _12883_/Q vssd1 vssd1 vccd1 vccd1 _10162_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput390 _11174_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10093_ _07886_/Y _10090_/X _08442_/Y _10047_/B vssd1 vssd1 vccd1 vccd1 _10093_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ _12890_/CLK _12803_/D _08355_/X vssd1 vssd1 vccd1 vccd1 _12803_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10995_ _11000_/D vssd1 vssd1 vccd1 vccd1 _10995_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12734_ _12749_/CLK _12734_/D _08617_/X vssd1 vssd1 vccd1 vccd1 _12734_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _13268_/CLK _12665_/D _08807_/X vssd1 vssd1 vccd1 vccd1 _12665_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _12970_/Q _12983_/Q _12601_/Q vssd1 vssd1 vccd1 vccd1 _11616_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _12939_/CLK _12596_/D vssd1 vssd1 vccd1 vccd1 _12596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11547_ _12804_/Q _09184_/A _11558_/S vssd1 vssd1 vccd1 vccd1 _11547_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11478_ _12921_/Q _10794_/B _11481_/S vssd1 vssd1 vccd1 vccd1 _11478_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13217_ _13217_/CLK _13217_/D _06622_/X vssd1 vssd1 vccd1 vccd1 _13217_/Q sky130_fd_sc_hd__dfrtp_1
X_10429_ _10429_/A _10429_/B _10429_/C vssd1 vssd1 vccd1 vccd1 _10433_/C sky130_fd_sc_hd__or3_4
XFILLER_98_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13148_ _13152_/CLK _13148_/D _07078_/X vssd1 vssd1 vccd1 vccd1 _13148_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13079_ _13081_/CLK _13079_/D _07292_/X vssd1 vssd1 vccd1 vccd1 _13079_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07640_ _12956_/Q _12954_/Q _07664_/A vssd1 vssd1 vccd1 vccd1 _07642_/B sky130_fd_sc_hd__or3_4
XFILLER_20_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07571_ _09982_/B _09441_/A _09435_/B vssd1 vssd1 vccd1 vccd1 _09439_/A sky130_fd_sc_hd__or3_4
XFILLER_20_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09310_ _12428_/Q _12427_/Q vssd1 vssd1 vccd1 vccd1 _09310_/X sky130_fd_sc_hd__or2_1
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06522_ _06522_/A vssd1 vssd1 vccd1 vccd1 _06522_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09241_ _12459_/Q _09231_/X _07568_/X _09233_/X vssd1 vssd1 vccd1 vccd1 _12459_/D
+ sky130_fd_sc_hd__a22o_1
X_06453_ _06458_/A _06458_/B vssd1 vssd1 vccd1 vccd1 _06453_/Y sky130_fd_sc_hd__nand2_1
XFILLER_142_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_90_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _13154_/CLK sky130_fd_sc_hd__clkbuf_16
X_09172_ _11621_/X _09163_/A _12496_/Q _09164_/A vssd1 vssd1 vccd1 vccd1 _12496_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06384_ _06382_/X _12220_/X _06375_/X _06383_/X vssd1 vssd1 vccd1 vccd1 _13247_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08123_ _12817_/Q vssd1 vssd1 vccd1 vccd1 _10439_/A sky130_fd_sc_hd__inv_2
XFILLER_107_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08054_ _08284_/A vssd1 vssd1 vccd1 vccd1 _08070_/A sky130_fd_sc_hd__buf_2
XFILLER_179_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07005_ _06457_/X _09524_/B _06459_/X _07004_/X vssd1 vssd1 vccd1 vccd1 _13173_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_1_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput107 la_data_in[46] vssd1 vssd1 vccd1 vccd1 input107/X sky130_fd_sc_hd__buf_1
Xinput118 la_data_in[56] vssd1 vssd1 vccd1 vccd1 input118/X sky130_fd_sc_hd__buf_1
X_08956_ _12468_/Q vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__inv_2
XFILLER_102_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput129 la_data_in[66] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_hd__buf_1
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07907_ _07967_/S vssd1 vssd1 vccd1 vccd1 _07918_/S sky130_fd_sc_hd__buf_2
XFILLER_5_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08887_ _08883_/X _06291_/Y _08878_/X _12634_/Q vssd1 vssd1 vccd1 vccd1 _12634_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07838_ _12905_/Q vssd1 vssd1 vccd1 vccd1 _10352_/B sky130_fd_sc_hd__inv_2
XFILLER_17_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07769_ _07769_/A vssd1 vssd1 vccd1 vccd1 _07769_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09508_ _13150_/Q _07737_/A _09507_/Y _09478_/X vssd1 vssd1 vccd1 vccd1 _09508_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_198_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10780_ _10779_/X _10731_/X _06389_/X _10732_/X _10733_/X vssd1 vssd1 vccd1 vccd1
+ _10780_/X sky130_fd_sc_hd__a221o_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09439_ _09439_/A vssd1 vssd1 vccd1 vccd1 _09440_/A sky130_fd_sc_hd__inv_2
XFILLER_13_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _12619_/CLK _12450_/D vssd1 vssd1 vccd1 vccd1 _12450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11401_ _10601_/Y _12408_/D _11404_/S vssd1 vssd1 vccd1 vccd1 _11401_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12381_ _12471_/CLK _12381_/D vssd1 vssd1 vccd1 vccd1 _12403_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_126_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11332_ vssd1 vssd1 vccd1 vccd1 _11332_/HI _11332_/LO sky130_fd_sc_hd__conb_1
XFILLER_126_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11263_ vssd1 vssd1 vccd1 vccd1 _11263_/HI _11263_/LO sky130_fd_sc_hd__conb_1
XFILLER_134_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13002_ _13004_/CLK _13002_/D vssd1 vssd1 vccd1 vccd1 _13002_/Q sky130_fd_sc_hd__dfxtp_1
X_10214_ _12663_/Q vssd1 vssd1 vccd1 vccd1 _10214_/Y sky130_fd_sc_hd__inv_2
X_11194_ vssd1 vssd1 vccd1 vccd1 _11194_/HI _11194_/LO sky130_fd_sc_hd__conb_1
XFILLER_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10145_ _12643_/Q vssd1 vssd1 vccd1 vccd1 _10145_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10076_ _12879_/Q vssd1 vssd1 vccd1 vccd1 _10076_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10978_ _10969_/Y _10970_/Y _10962_/Y _10963_/Y vssd1 vssd1 vccd1 vccd1 _10978_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ _12717_/CLK _12717_/D _08661_/X vssd1 vssd1 vccd1 vccd1 _12717_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ _12653_/CLK _12648_/D _08848_/X vssd1 vssd1 vccd1 vccd1 _12648_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12579_ _12992_/CLK _12579_/D vssd1 vssd1 vccd1 vccd1 _12579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08810_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08810_/X sky130_fd_sc_hd__clkbuf_1
X_09790_ _09790_/A vssd1 vssd1 vccd1 vccd1 _09790_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08741_ _08741_/A vssd1 vssd1 vccd1 vccd1 _08764_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08672_ _11847_/X _08670_/X _12713_/Q _08671_/X vssd1 vssd1 vccd1 vccd1 _12713_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07623_ _12962_/Q vssd1 vssd1 vccd1 vccd1 _07661_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07554_ _07775_/A vssd1 vssd1 vccd1 vccd1 _09002_/A sky130_fd_sc_hd__buf_2
XFILLER_22_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06505_ _06440_/X _06503_/Y _06489_/X _06504_/Y vssd1 vssd1 vccd1 vccd1 _13228_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07485_ _07489_/A vssd1 vssd1 vccd1 vccd1 _07485_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09224_ _12468_/Q _11803_/X _09224_/S vssd1 vssd1 vccd1 vccd1 _12468_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06436_ _06887_/A vssd1 vssd1 vccd1 vccd1 _06436_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_107_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09155_ _09155_/A vssd1 vssd1 vccd1 vccd1 _09164_/A sky130_fd_sc_hd__inv_2
X_06367_ _06370_/A vssd1 vssd1 vccd1 vccd1 _06367_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08106_ _12808_/Q vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__inv_2
XFILLER_108_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09086_ _12542_/Q _09079_/Y _09179_/B _09083_/X vssd1 vssd1 vccd1 vccd1 _12542_/D
+ sky130_fd_sc_hd__o22a_1
X_06298_ _06087_/Y _06088_/Y _06091_/B _06179_/Y vssd1 vssd1 vccd1 vccd1 _06298_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08037_ _12871_/Q _08024_/X _07993_/X _08026_/X vssd1 vssd1 vccd1 vccd1 _12871_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09988_ _09980_/Y _10163_/A _09679_/Y _10166_/A _09987_/X vssd1 vssd1 vccd1 vccd1
+ _09988_/X sky130_fd_sc_hd__o221a_1
XFILLER_104_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08939_ _12435_/Q _12121_/S vssd1 vssd1 vccd1 vccd1 _08940_/B sky130_fd_sc_hd__and2b_1
XFILLER_88_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11950_ _09809_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11950_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10901_ _10900_/A _10900_/B _10900_/Y vssd1 vssd1 vccd1 vccd1 _10903_/A sky130_fd_sc_hd__a21oi_2
XFILLER_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11881_ _11051_/Y _10731_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _11881_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10832_ _10824_/Y _10825_/Y _10827_/Y _10828_/Y vssd1 vssd1 vccd1 vccd1 _10832_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_199_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10763_ _10763_/A vssd1 vssd1 vccd1 vccd1 _10763_/X sky130_fd_sc_hd__buf_2
XFILLER_125_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12502_ _13244_/CLK _12502_/D vssd1 vssd1 vccd1 vccd1 _12502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10694_ _06407_/X _10691_/A _10691_/B _10693_/X _10701_/A vssd1 vssd1 vccd1 vccd1
+ _10694_/X sky130_fd_sc_hd__a32o_1
XFILLER_201_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12433_ _12480_/CLK _12433_/D vssd1 vssd1 vccd1 vccd1 _12433_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ _12620_/CLK _12364_/D vssd1 vssd1 vccd1 vccd1 _12364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11315_ vssd1 vssd1 vccd1 vccd1 _11315_/HI _11315_/LO sky130_fd_sc_hd__conb_1
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12295_ _12558_/CLK _12295_/D vssd1 vssd1 vccd1 vccd1 _12295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11246_ vssd1 vssd1 vccd1 vccd1 _11246_/HI _11246_/LO sky130_fd_sc_hd__conb_1
XFILLER_45_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11177_ vssd1 vssd1 vccd1 vccd1 _11177_/HI _11177_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10128_ _10128_/A _10128_/B _10128_/C _10128_/D vssd1 vssd1 vccd1 vccd1 _10128_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_110_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10059_ _12639_/Q vssd1 vssd1 vccd1 vccd1 _10059_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12422_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07270_ _07280_/A vssd1 vssd1 vccd1 vccd1 _07270_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06221_ _06245_/A vssd1 vssd1 vccd1 vccd1 _06221_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06152_ _12746_/Q _12714_/Q _12745_/Q _12713_/Q vssd1 vssd1 vccd1 vccd1 _06152_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06083_ _12697_/Q vssd1 vssd1 vccd1 vccd1 _06083_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09911_ _09909_/Y _09897_/X _06323_/A _09892_/X _09910_/X vssd1 vssd1 vccd1 vccd1
+ _09911_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_99_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09842_ _09842_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _09842_/X sky130_fd_sc_hd__or2_1
XFILLER_99_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09773_ _09717_/B _09770_/X _09717_/A _09770_/X _09829_/A vssd1 vssd1 vccd1 vccd1
+ _09785_/A sky130_fd_sc_hd__o221a_1
X_06985_ _07006_/A vssd1 vssd1 vccd1 vccd1 _06985_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08724_ _11826_/X _08715_/X _12692_/Q _08716_/X vssd1 vssd1 vccd1 vccd1 _12692_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _08686_/A vssd1 vssd1 vccd1 vccd1 _08655_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _07599_/Y _07600_/B _07605_/Y _09002_/A vssd1 vssd1 vccd1 vccd1 _12975_/D
+ sky130_fd_sc_hd__a31oi_1
XPHY_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _11955_/X _08575_/X _12746_/Q _08578_/X vssd1 vssd1 vccd1 vccd1 _12746_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07537_ _13000_/Q _07531_/X _07536_/X _07532_/X _09023_/A vssd1 vssd1 vccd1 vccd1
+ _13000_/D sky130_fd_sc_hd__o221a_1
XPHY_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07468_ _11460_/X _07459_/X _13019_/Q _07460_/X vssd1 vssd1 vccd1 vccd1 _13019_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09207_ _09215_/A vssd1 vssd1 vccd1 vccd1 _09207_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06419_ _06886_/A vssd1 vssd1 vccd1 vccd1 _06769_/A sky130_fd_sc_hd__buf_2
XFILLER_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07399_ _11419_/X _07368_/A _13043_/Q _07369_/A vssd1 vssd1 vccd1 vccd1 _13043_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09138_ _12499_/Q _09138_/B vssd1 vssd1 vccd1 vccd1 _09139_/B sky130_fd_sc_hd__or2_1
XFILLER_108_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09069_ _11147_/A vssd1 vssd1 vccd1 vccd1 _09069_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_191_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11100_ _11100_/A vssd1 vssd1 vccd1 vccd1 _11100_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12080_ _12447_/Q _10683_/X _12090_/S vssd1 vssd1 vccd1 vccd1 _12080_/X sky130_fd_sc_hd__mux2_1
X_11031_ _11031_/A vssd1 vssd1 vccd1 vccd1 _12614_/D sky130_fd_sc_hd__inv_2
XFILLER_134_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12982_ _13001_/CLK _12982_/D vssd1 vssd1 vccd1 vccd1 _12982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11933_ _09543_/X _12794_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11933_/X sky130_fd_sc_hd__mux2_2
XFILLER_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11864_ _10129_/Y _12317_/Q _12312_/Q vssd1 vssd1 vccd1 vccd1 _11864_/X sky130_fd_sc_hd__mux2_2
XPHY_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10815_ _12326_/Q vssd1 vssd1 vccd1 vccd1 _10815_/Y sky130_fd_sc_hd__inv_2
XPHY_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11795_ _12060_/X _12483_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11795_/X sky130_fd_sc_hd__mux2_1
XPHY_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10746_ _11054_/A vssd1 vssd1 vccd1 vccd1 _10746_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_147_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12550_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10677_ _12439_/Q _09315_/A _12439_/Q _09315_/A vssd1 vssd1 vccd1 vccd1 _10677_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12416_ _12467_/CLK _12416_/D vssd1 vssd1 vccd1 vccd1 _12416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12347_ _12541_/CLK _12347_/D vssd1 vssd1 vccd1 vccd1 _12347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12278_ _10262_/X _12904_/Q _11874_/X _10260_/Y _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12294_/D sky130_fd_sc_hd__mux4_2
XFILLER_107_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11229_ vssd1 vssd1 vccd1 vccd1 _11229_/HI _11229_/LO sky130_fd_sc_hd__conb_1
XFILLER_95_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06770_ _06757_/X _06761_/X _06762_/X vssd1 vssd1 vccd1 vccd1 _06770_/X sky130_fd_sc_hd__a21bo_1
XFILLER_83_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput290 la_oenb[96] vssd1 vssd1 vccd1 vccd1 input290/X sky130_fd_sc_hd__buf_1
XFILLER_36_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08440_ _13046_/Q vssd1 vssd1 vccd1 vccd1 _08440_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08371_ _12798_/Q _08358_/X _07993_/X _08360_/X vssd1 vssd1 vccd1 vccd1 _12798_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07322_ _07384_/A vssd1 vssd1 vccd1 vccd1 _07385_/A sky130_fd_sc_hd__inv_2
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07253_ _07253_/A vssd1 vssd1 vccd1 vccd1 _07266_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_192_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06204_ _06030_/A _06198_/X _06030_/A _06198_/X vssd1 vssd1 vccd1 vccd1 _06204_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_9_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07184_ _11519_/X _07176_/X _13118_/Q _07177_/X vssd1 vssd1 vccd1 vccd1 _13118_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06135_ _12738_/Q _12706_/Q _12737_/Q _12705_/Q vssd1 vssd1 vccd1 vccd1 _06135_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06066_ _12702_/Q vssd1 vssd1 vccd1 vccd1 _06067_/B sky130_fd_sc_hd__inv_2
XFILLER_160_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09825_ _09825_/A vssd1 vssd1 vccd1 vccd1 _09825_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09756_ _09738_/Y _06677_/Y _06659_/Y _09740_/Y vssd1 vssd1 vccd1 vccd1 _09756_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06968_ _06961_/Y _06966_/Y _06971_/A vssd1 vssd1 vccd1 vccd1 _06977_/A sky130_fd_sc_hd__o21ba_1
XFILLER_101_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08707_ _11833_/X _08700_/X _12699_/Q _08701_/X vssd1 vssd1 vccd1 vccd1 _12699_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09687_ _06792_/Y _06796_/Y _09665_/Y _09666_/Y vssd1 vssd1 vccd1 vccd1 _09687_/X
+ sky130_fd_sc_hd__o22a_4
X_06899_ _12024_/X _12020_/X _06898_/X vssd1 vssd1 vccd1 vccd1 _06899_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _08638_/A vssd1 vssd1 vccd1 vccd1 _08638_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _08569_/A vssd1 vssd1 vccd1 vccd1 _08569_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ _12407_/D _12408_/D _10603_/B vssd1 vssd1 vccd1 vccd1 _10600_/X sky130_fd_sc_hd__o21a_1
XPHY_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ _10408_/X _09185_/D _11610_/S vssd1 vssd1 vccd1 vccd1 _11580_/X sky130_fd_sc_hd__mux2_1
XPHY_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10531_ _12321_/Q _09327_/B _10608_/A _12363_/Q vssd1 vssd1 vccd1 vccd1 _10532_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13250_ _13252_/CLK _13250_/D _06370_/X vssd1 vssd1 vccd1 vccd1 _13250_/Q sky130_fd_sc_hd__dfrtp_2
X_10462_ _10462_/A vssd1 vssd1 vccd1 vccd1 _10462_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12201_ _11132_/X _10776_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12201_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13181_ _13183_/CLK _13181_/D _06942_/X vssd1 vssd1 vccd1 vccd1 _13181_/Q sky130_fd_sc_hd__dfrtp_1
X_10393_ _10393_/A _10393_/B vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__or2_4
XFILLER_2_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12132_ _10707_/Y _06468_/A _12766_/Q vssd1 vssd1 vccd1 vccd1 _12132_/X sky130_fd_sc_hd__mux2_2
XFILLER_2_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12063_ _12440_/Q _12062_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12063_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11014_ _11014_/A _11014_/B _11014_/C _11014_/D vssd1 vssd1 vccd1 vccd1 _11018_/C
+ sky130_fd_sc_hd__nor4_2
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12965_ _12976_/CLK _12965_/D vssd1 vssd1 vccd1 vccd1 _12965_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11916_ _10657_/X _09317_/X _11916_/S vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12896_ _12166_/X _12896_/D _07959_/X vssd1 vssd1 vccd1 vccd1 _12896_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _09958_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11777_/X _12125_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12434_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10729_ _13253_/Q _06425_/A _10730_/A _10717_/X _06430_/A vssd1 vssd1 vccd1 vccd1
+ _11146_/A sky130_fd_sc_hd__o221a_1
XFILLER_119_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07940_ _12904_/Q _11493_/X _07946_/S vssd1 vssd1 vccd1 vccd1 _12904_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12985_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07871_ _12922_/Q vssd1 vssd1 vccd1 vccd1 _10395_/A sky130_fd_sc_hd__clkinv_4
XFILLER_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09610_ _09574_/B _09632_/A _09558_/B _09608_/Y _09609_/X vssd1 vssd1 vccd1 vccd1
+ _09611_/B sky130_fd_sc_hd__o311a_1
X_06822_ _13196_/Q vssd1 vssd1 vccd1 vccd1 _06822_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09541_ _09528_/A _09530_/X _09540_/Y vssd1 vssd1 vccd1 vccd1 _09541_/Y sky130_fd_sc_hd__o21ai_1
X_06753_ _12014_/X _06728_/X _12014_/X _06728_/X vssd1 vssd1 vccd1 vccd1 _06754_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09472_ _13164_/Q vssd1 vssd1 vccd1 vccd1 _09482_/A sky130_fd_sc_hd__inv_2
X_06684_ _06658_/X _06677_/Y _06608_/X _06683_/X vssd1 vssd1 vccd1 vccd1 _13211_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ _08433_/A vssd1 vssd1 vccd1 vccd1 _08423_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ _08372_/A vssd1 vssd1 vccd1 vccd1 _08370_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07305_ _13076_/Q _07285_/X _07304_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _13076_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08285_ _08296_/A vssd1 vssd1 vccd1 vccd1 _08285_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07236_ _07236_/A vssd1 vssd1 vccd1 vccd1 _07236_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07167_ _07167_/A vssd1 vssd1 vccd1 vccd1 _07167_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06118_ _12687_/Q vssd1 vssd1 vccd1 vccd1 _06118_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07098_ _07098_/A _07098_/B vssd1 vssd1 vccd1 vccd1 _09041_/B sky130_fd_sc_hd__or2_1
Xoutput550 _11295_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__clkbuf_2
Xoutput561 _11305_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__clkbuf_2
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput572 _11315_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__clkbuf_2
X_06049_ _12739_/Q _12707_/Q _06047_/Y _06048_/Y vssd1 vssd1 vccd1 vccd1 _06051_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput583 _12556_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput594 _12566_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09808_ _09823_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09808_/X sky130_fd_sc_hd__or2_1
XFILLER_47_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09739_ _13212_/Q _13211_/Q _09738_/Y _06677_/Y vssd1 vssd1 vccd1 vccd1 _09740_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _13256_/CLK _12750_/D _08560_/X vssd1 vssd1 vccd1 vccd1 _12750_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11887_/X _09180_/B _11703_/S vssd1 vssd1 vccd1 vccd1 _11701_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12681_ _12682_/CLK _12681_/D _08755_/X vssd1 vssd1 vccd1 vccd1 _12681_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _10502_/X _12931_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11632_/X sky130_fd_sc_hd__mux2_1
XPHY_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ _12820_/Q _09179_/B _11569_/S vssd1 vssd1 vccd1 vccd1 _11563_/X sky130_fd_sc_hd__mux2_1
XPHY_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10514_ _12588_/Q _07762_/B _07763_/B vssd1 vssd1 vccd1 vccd1 _10514_/X sky130_fd_sc_hd__a21bo_1
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11494_ _10351_/X _09244_/A _11501_/S vssd1 vssd1 vccd1 vccd1 _11494_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13233_ _13237_/CLK _13233_/D _06461_/X vssd1 vssd1 vccd1 vccd1 _13233_/Q sky130_fd_sc_hd__dfrtp_1
X_10445_ _10455_/D vssd1 vssd1 vccd1 vccd1 _10447_/B sky130_fd_sc_hd__inv_2
XFILLER_124_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13164_ _13254_/CLK _13164_/D _07029_/X vssd1 vssd1 vccd1 vccd1 _13164_/Q sky130_fd_sc_hd__dfrtp_4
X_10376_ _12914_/Q _12913_/Q _10376_/C vssd1 vssd1 vccd1 vccd1 _10377_/A sky130_fd_sc_hd__and3_1
X_12115_ _12114_/X _12433_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12115_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13095_ _12167_/X _13095_/D _07247_/X vssd1 vssd1 vccd1 vccd1 _13095_/Q sky130_fd_sc_hd__dfrtp_4
X_12046_ _10719_/X _11129_/A _12193_/S vssd1 vssd1 vccd1 vccd1 _12046_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12948_ _12951_/CLK _12948_/D vssd1 vssd1 vccd1 vccd1 _12948_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_162_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12535_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ _12880_/CLK _12879_/D _08014_/X vssd1 vssd1 vccd1 vccd1 _12879_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08070_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07021_ _06886_/X _07020_/X _06887_/X _13168_/Q vssd1 vssd1 vccd1 vccd1 _13168_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_161_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08972_ _09067_/A vssd1 vssd1 vccd1 vccd1 _08972_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07923_ _07931_/A vssd1 vssd1 vccd1 vccd1 _07923_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07854_ _12912_/Q vssd1 vssd1 vccd1 vccd1 _10367_/A sky130_fd_sc_hd__inv_2
XFILLER_29_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06805_ _06719_/X _06800_/X _06804_/Y _06480_/X _13197_/Q vssd1 vssd1 vccd1 vccd1
+ _13197_/D sky130_fd_sc_hd__a32o_1
X_07785_ _07560_/X _07780_/X _12930_/Q _07781_/X _07775_/X vssd1 vssd1 vccd1 vccd1
+ _12930_/D sky130_fd_sc_hd__a221o_1
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09524_ _09524_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09524_/Y sky130_fd_sc_hd__nor2_2
X_06736_ _06630_/X _06730_/X _06734_/X _06646_/X _06735_/Y vssd1 vssd1 vccd1 vccd1
+ _06737_/A sky130_fd_sc_hd__a32o_1
XFILLER_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _12981_/Q _09436_/A _12997_/Q _09451_/X vssd1 vssd1 vccd1 vccd1 _09455_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06667_ _12048_/X _12047_/X _12048_/X _12047_/X vssd1 vssd1 vccd1 vccd1 _06667_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ _12786_/Q _08401_/X _07980_/X _08403_/X vssd1 vssd1 vccd1 vccd1 _12786_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09386_ _12453_/Q _09384_/Y _12458_/Q _09385_/Y vssd1 vssd1 vccd1 vccd1 _09386_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06598_ _06598_/A _06598_/B vssd1 vssd1 vccd1 vccd1 _06598_/Y sky130_fd_sc_hd__nor2_2
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08337_ _08337_/A vssd1 vssd1 vccd1 vccd1 _08349_/S sky130_fd_sc_hd__buf_2
XFILLER_138_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08268_ _08282_/A vssd1 vssd1 vccd1 vccd1 _08268_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07219_ _07249_/A vssd1 vssd1 vccd1 vccd1 _07219_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_180_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08199_ _13089_/Q vssd1 vssd1 vccd1 vccd1 _08199_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10230_ _13091_/Q _10228_/X _13123_/Q _10229_/X vssd1 vssd1 vccd1 vccd1 _10230_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10161_ _12867_/Q vssd1 vssd1 vccd1 vccd1 _10161_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput380 _11165_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput391 _11175_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10092_ _08194_/Y _10070_/X _10091_/X vssd1 vssd1 vccd1 vccd1 _10092_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_120_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12802_ _12802_/CLK _12802_/D _08362_/X vssd1 vssd1 vccd1 vccd1 _12802_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_90_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10994_ _12541_/Q _12353_/Q _10993_/X vssd1 vssd1 vccd1 vccd1 _11000_/D sky130_fd_sc_hd__a21bo_1
XFILLER_90_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12733_ _12749_/CLK _12733_/D _08619_/X vssd1 vssd1 vccd1 vccd1 _12733_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12664_/CLK _12664_/D _08810_/X vssd1 vssd1 vccd1 vccd1 _12664_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _12969_/Q _12982_/Q _12601_/Q vssd1 vssd1 vccd1 vccd1 _11615_/X sky130_fd_sc_hd__mux2_1
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ _12973_/CLK _12595_/D vssd1 vssd1 vccd1 vccd1 _12595_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ _12835_/Q _10793_/A _11546_/S vssd1 vssd1 vccd1 vccd1 _11546_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11477_ _12920_/Q _10794_/C _11481_/S vssd1 vssd1 vccd1 vccd1 _11477_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13216_ _13217_/CLK _13216_/D _06624_/X vssd1 vssd1 vccd1 vccd1 _13216_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10428_ _10429_/B _10429_/C _10429_/A vssd1 vssd1 vccd1 vccd1 _10431_/A sky130_fd_sc_hd__o21a_1
XFILLER_100_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13147_ _13152_/CLK _13147_/D _07081_/X vssd1 vssd1 vccd1 vccd1 _13147_/Q sky130_fd_sc_hd__dfrtp_2
X_10359_ _10357_/B _10357_/C _10357_/A vssd1 vssd1 vccd1 vccd1 _10360_/C sky130_fd_sc_hd__o21a_1
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13078_ _13081_/CLK _13078_/D _07295_/X vssd1 vssd1 vccd1 vccd1 _13078_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12029_ _11121_/X _11114_/X _12193_/S vssd1 vssd1 vccd1 vccd1 _12029_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07570_ _07568_/X _07552_/A _12986_/Q _07553_/A _07569_/X vssd1 vssd1 vccd1 vccd1
+ _12986_/D sky130_fd_sc_hd__a221o_1
XFILLER_20_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06521_ _06507_/X _06508_/Y _06489_/X _06520_/Y vssd1 vssd1 vccd1 vccd1 _13227_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09240_ _12460_/Q _09231_/X _07566_/X _09233_/X vssd1 vssd1 vccd1 vccd1 _12460_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06452_ _06444_/A _06444_/B _06451_/Y _06444_/Y _06451_/A vssd1 vssd1 vccd1 vccd1
+ _06458_/B sky130_fd_sc_hd__o32a_1
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09171_ _11622_/X _09163_/A _12497_/Q _09164_/A vssd1 vssd1 vccd1 vccd1 _12497_/D
+ sky130_fd_sc_hd__a22o_1
X_06383_ _13247_/Q vssd1 vssd1 vccd1 vccd1 _06383_/X sky130_fd_sc_hd__buf_2
XFILLER_193_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08122_ _12835_/Q vssd1 vssd1 vccd1 vccd1 _08122_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08053_ _08657_/A vssd1 vssd1 vccd1 vccd1 _08284_/A sky130_fd_sc_hd__buf_2
X_07004_ _06999_/Y _11853_/X _07003_/Y vssd1 vssd1 vccd1 vccd1 _07004_/X sky130_fd_sc_hd__o21a_1
XFILLER_116_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08955_ _10627_/A vssd1 vssd1 vccd1 vccd1 _12103_/S sky130_fd_sc_hd__clkinv_4
Xinput108 la_data_in[47] vssd1 vssd1 vccd1 vccd1 input108/X sky130_fd_sc_hd__buf_1
Xinput119 la_data_in[57] vssd1 vssd1 vccd1 vccd1 input119/X sky130_fd_sc_hd__buf_1
XFILLER_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07906_ _07917_/A vssd1 vssd1 vccd1 vccd1 _07906_/X sky130_fd_sc_hd__clkbuf_1
X_08886_ _08897_/A vssd1 vssd1 vccd1 vccd1 _08886_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07837_ _12913_/Q vssd1 vssd1 vccd1 vccd1 _10373_/A sky130_fd_sc_hd__inv_2
XFILLER_45_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07768_ _07768_/A vssd1 vssd1 vccd1 vccd1 _11648_/S sky130_fd_sc_hd__buf_8
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09507_ _12864_/Q vssd1 vssd1 vccd1 vccd1 _09507_/Y sky130_fd_sc_hd__inv_2
X_06719_ _06887_/A vssd1 vssd1 vccd1 vccd1 _06719_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_197_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07699_ _12961_/Q _07694_/X _12960_/Q _07698_/X _07695_/X vssd1 vssd1 vccd1 vccd1
+ _12961_/D sky130_fd_sc_hd__o221a_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09438_/A vssd1 vssd1 vccd1 vccd1 _09438_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_198_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09369_ _12454_/Q _09367_/Y _12546_/Q _09368_/Y vssd1 vssd1 vccd1 vccd1 _09369_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11400_ _10604_/X _12409_/D _11403_/S vssd1 vssd1 vccd1 vccd1 _11400_/X sky130_fd_sc_hd__mux2_1
X_12380_ _13008_/CLK _12380_/D vssd1 vssd1 vccd1 vccd1 _12402_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_166_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11331_ vssd1 vssd1 vccd1 vccd1 _11331_/HI _11331_/LO sky130_fd_sc_hd__conb_1
XFILLER_181_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11262_ vssd1 vssd1 vccd1 vccd1 _11262_/HI _11262_/LO sky130_fd_sc_hd__conb_1
X_13001_ _13001_/CLK _13001_/D vssd1 vssd1 vccd1 vccd1 _13001_/Q sky130_fd_sc_hd__dfxtp_2
X_10213_ _07820_/Y _10151_/X _10212_/X vssd1 vssd1 vccd1 vccd1 _10213_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11193_ vssd1 vssd1 vccd1 vccd1 _11193_/HI _11193_/LO sky130_fd_sc_hd__conb_1
XFILLER_161_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10144_ _13152_/Q vssd1 vssd1 vccd1 vccd1 _10144_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10075_ _12624_/Q vssd1 vssd1 vccd1 vccd1 _10075_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10977_ _10977_/A _10977_/B _10977_/C _10977_/D vssd1 vssd1 vccd1 vccd1 _10980_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12716_ _12716_/CLK _12716_/D _08663_/X vssd1 vssd1 vccd1 vccd1 _12716_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12647_ _12753_/CLK _12647_/D _08851_/X vssd1 vssd1 vccd1 vccd1 _12647_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_175_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12578_ _12976_/CLK _12578_/D vssd1 vssd1 vccd1 vccd1 _12578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11529_ _12818_/Q _09243_/A _11533_/S vssd1 vssd1 vccd1 vccd1 _11529_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08740_ _08740_/A _08811_/A vssd1 vssd1 vccd1 vccd1 _08741_/A sky130_fd_sc_hd__or2_1
XFILLER_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08671_ _08686_/A vssd1 vssd1 vccd1 vccd1 _08671_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07622_ _12946_/Q vssd1 vssd1 vccd1 vccd1 _07678_/B sky130_fd_sc_hd__inv_2
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07553_ _07553_/A vssd1 vssd1 vccd1 vccd1 _07553_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06504_ _06500_/A _06500_/B _06500_/Y vssd1 vssd1 vccd1 vccd1 _06504_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07484_ _11454_/X _07474_/X _13013_/Q _07475_/X vssd1 vssd1 vccd1 vccd1 _13013_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09223_ _12449_/Q _09304_/B vssd1 vssd1 vccd1 vccd1 _09224_/S sky130_fd_sc_hd__or2b_1
XFILLER_195_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06435_ _06841_/A vssd1 vssd1 vccd1 vccd1 _06435_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_146_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09154_ _09163_/A vssd1 vssd1 vccd1 vccd1 _09154_/X sky130_fd_sc_hd__clkbuf_2
X_06366_ _06361_/X _12230_/X _06358_/X _06365_/X vssd1 vssd1 vccd1 vccd1 _13252_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08105_ _13118_/Q vssd1 vssd1 vccd1 vccd1 _08105_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09085_ _12543_/Q _09079_/Y _09179_/A _09083_/X vssd1 vssd1 vccd1 vccd1 _12543_/D
+ sky130_fd_sc_hd__o22a_1
X_06297_ _06313_/A vssd1 vssd1 vccd1 vccd1 _06297_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08036_ _08036_/A vssd1 vssd1 vccd1 vccd1 _08036_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 la_data_in[30] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__buf_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09987_ _09983_/Y _10165_/A _09985_/Y _10168_/A vssd1 vssd1 vccd1 vccd1 _09987_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08938_ _12433_/Q _12434_/Q vssd1 vssd1 vccd1 vccd1 _12121_/S sky130_fd_sc_hd__nor2_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08869_ _08882_/A vssd1 vssd1 vccd1 vccd1 _08869_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10900_ _10900_/A _10900_/B vssd1 vssd1 vccd1 vccd1 _10900_/Y sky130_fd_sc_hd__nor2_2
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11880_ _11099_/A _10708_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _11880_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10831_ _12517_/Q _12329_/Q _10830_/X vssd1 vssd1 vccd1 vccd1 _10831_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_199_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10762_ _10758_/X _10759_/X _06376_/X _10760_/X _10761_/X vssd1 vssd1 vccd1 vccd1
+ _10762_/X sky130_fd_sc_hd__a221o_1
XFILLER_197_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12501_ _13243_/CLK _12501_/D vssd1 vssd1 vccd1 vccd1 _12501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10693_ _10693_/A vssd1 vssd1 vccd1 vccd1 _10693_/X sky130_fd_sc_hd__buf_2
XFILLER_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12432_ _12480_/CLK _12432_/D vssd1 vssd1 vccd1 vccd1 _12432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ _12376_/CLK _12363_/D vssd1 vssd1 vccd1 vccd1 _12363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11314_ vssd1 vssd1 vccd1 vccd1 _11314_/HI _11314_/LO sky130_fd_sc_hd__conb_1
XFILLER_153_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12294_ _12296_/CLK _12294_/D vssd1 vssd1 vccd1 vccd1 _12294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11245_ vssd1 vssd1 vccd1 vccd1 _11245_/HI _11245_/LO sky130_fd_sc_hd__conb_1
XFILLER_106_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11176_ vssd1 vssd1 vccd1 vccd1 _11176_/HI _11176_/LO sky130_fd_sc_hd__conb_1
XFILLER_110_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10127_ _10123_/Y _09999_/A _10124_/Y _10141_/A _10126_/X vssd1 vssd1 vccd1 vccd1
+ _10128_/D sky130_fd_sc_hd__o221a_1
XFILLER_95_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10058_ _10056_/Y _10018_/X _10057_/Y _10020_/X vssd1 vssd1 vccd1 vccd1 _10068_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_69_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12976_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_177_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06220_ _08996_/D vssd1 vssd1 vccd1 vccd1 _06245_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06151_ _06185_/A _06151_/B vssd1 vssd1 vccd1 vccd1 _06151_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06082_ _12729_/Q vssd1 vssd1 vccd1 vccd1 _06082_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09910_ _12883_/Q _09910_/B vssd1 vssd1 vccd1 vccd1 _09910_/X sky130_fd_sc_hd__or2_1
XFILLER_98_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09841_ _09842_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _09841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09772_ _09749_/Y _09803_/A _09771_/Y vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__o21a_1
XFILLER_86_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06984_ _06528_/X _06965_/X _06983_/Y _06841_/X _13176_/Q vssd1 vssd1 vccd1 vccd1
+ _13176_/D sky130_fd_sc_hd__a32o_1
XFILLER_112_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08723_ _08729_/A vssd1 vssd1 vccd1 vccd1 _08723_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08654_ _08685_/A vssd1 vssd1 vccd1 vccd1 _08654_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07605_ _12974_/Q _07610_/A _12975_/Q vssd1 vssd1 vccd1 vccd1 _07605_/Y sky130_fd_sc_hd__o21ai_1
XPHY_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08585_ _08591_/A vssd1 vssd1 vccd1 vccd1 _08585_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07536_ _09184_/B vssd1 vssd1 vccd1 vccd1 _07536_/X sky130_fd_sc_hd__buf_4
XPHY_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07467_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07467_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09206_ _12481_/Q _09199_/X _09244_/A _09200_/X vssd1 vssd1 vccd1 vccd1 _12481_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06418_ _12621_/Q vssd1 vssd1 vccd1 vccd1 _06886_/A sky130_fd_sc_hd__inv_2
XFILLER_195_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07398_ _07408_/A vssd1 vssd1 vccd1 vccd1 _07398_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_124_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09137_ _12498_/Q _09137_/B vssd1 vssd1 vccd1 vccd1 _09138_/B sky130_fd_sc_hd__or2_1
XFILLER_33_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06349_ _06370_/A vssd1 vssd1 vccd1 vccd1 _06349_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09068_ _11147_/A vssd1 vssd1 vccd1 vccd1 _09068_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08019_ _12877_/Q _07996_/A _07313_/X _07998_/A vssd1 vssd1 vccd1 vccd1 _12877_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11030_ _12312_/Q _11030_/B vssd1 vssd1 vccd1 vccd1 _12312_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12981_ _13001_/CLK _12981_/D vssd1 vssd1 vccd1 vccd1 _12981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11932_ _09534_/Y _12793_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11932_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11863_ _10131_/X _12808_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _12514_/Q vssd1 vssd1 vccd1 vccd1 _10814_/Y sky130_fd_sc_hd__inv_2
XPHY_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _11793_/X _12143_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12438_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10745_ _10745_/A vssd1 vssd1 vccd1 vccd1 _11054_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_186_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10676_ _12437_/Q _12438_/Q vssd1 vssd1 vccd1 vccd1 _10676_/X sky130_fd_sc_hd__and2_1
XFILLER_139_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12415_ _12415_/CLK _12415_/D vssd1 vssd1 vccd1 vccd1 _12415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12346_ _12529_/CLK _12346_/D vssd1 vssd1 vccd1 vccd1 _12346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_116_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 _12717_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12277_ _10247_/X _12903_/Q _11873_/X _10245_/Y _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12293_/D sky130_fd_sc_hd__mux4_2
X_11228_ vssd1 vssd1 vccd1 vccd1 _11228_/HI _11228_/LO sky130_fd_sc_hd__conb_1
XFILLER_49_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ vssd1 vssd1 vccd1 vccd1 _11159_/HI _11159_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput280 la_oenb[87] vssd1 vssd1 vccd1 vccd1 input280/X sky130_fd_sc_hd__buf_1
Xinput291 la_oenb[97] vssd1 vssd1 vccd1 vccd1 input291/X sky130_fd_sc_hd__buf_1
XFILLER_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08370_ _08370_/A vssd1 vssd1 vccd1 vccd1 _08370_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07321_ _07368_/A vssd1 vssd1 vccd1 vccd1 _07321_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07252_ _11559_/X _07248_/X _13094_/Q _07249_/X vssd1 vssd1 vccd1 vccd1 _13094_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06203_ _13282_/Q vssd1 vssd1 vccd1 vccd1 _06203_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07183_ _07183_/A vssd1 vssd1 vccd1 vccd1 _07183_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06134_ _06134_/A vssd1 vssd1 vccd1 vccd1 _06134_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06065_ _12734_/Q vssd1 vssd1 vccd1 vccd1 _06067_/A sky130_fd_sc_hd__inv_2
XFILLER_28_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09824_ _09824_/A _09848_/A vssd1 vssd1 vccd1 vccd1 _09868_/C sky130_fd_sc_hd__or2_1
XFILLER_24_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09755_ _13217_/Q vssd1 vssd1 vccd1 vccd1 _09755_/Y sky130_fd_sc_hd__inv_2
X_06967_ _06961_/A _06961_/B _06961_/Y _06966_/Y vssd1 vssd1 vccd1 vccd1 _06971_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08706_ _08714_/A vssd1 vssd1 vccd1 vccd1 _08706_/X sky130_fd_sc_hd__clkbuf_1
X_09686_ _09686_/A vssd1 vssd1 vccd1 vccd1 _09686_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06898_ _12017_/X _06898_/B vssd1 vssd1 vccd1 vccd1 _06898_/X sky130_fd_sc_hd__or2_1
X_08637_ _11935_/X _08624_/X _12726_/Q _08625_/X vssd1 vssd1 vccd1 vccd1 _12726_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _08561_/Y _08565_/X _08552_/B _08567_/X vssd1 vssd1 vccd1 vccd1 _12750_/D
+ sky130_fd_sc_hd__o22ai_1
XPHY_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07519_ _13001_/Q _07519_/B vssd1 vssd1 vccd1 vccd1 _07520_/A sky130_fd_sc_hd__nand2_2
XPHY_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08499_ _12945_/Q vssd1 vssd1 vccd1 vccd1 _08499_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10530_ _12321_/Q vssd1 vssd1 vccd1 vccd1 _10608_/A sky130_fd_sc_hd__inv_2
XPHY_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10461_ _12824_/Q _10463_/C _10459_/X _10462_/A vssd1 vssd1 vccd1 vccd1 _10461_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12200_ _11131_/X _10775_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _12200_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ _13190_/CLK _13180_/D _06952_/X vssd1 vssd1 vccd1 vccd1 _13180_/Q sky130_fd_sc_hd__dfrtp_4
X_10392_ _10390_/A _10390_/B _10387_/A _10391_/Y vssd1 vssd1 vccd1 vccd1 _10392_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_108_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12131_ _10715_/Y _10714_/Y _12770_/Q vssd1 vssd1 vccd1 vccd1 _12131_/X sky130_fd_sc_hd__mux2_2
XFILLER_190_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12062_ _12061_/X _12440_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12062_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_11013_ _11013_/A _11013_/B vssd1 vssd1 vccd1 vccd1 _11014_/C sky130_fd_sc_hd__or2_1
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12964_ _12976_/CLK _12964_/D vssd1 vssd1 vccd1 vccd1 _12964_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11915_ _11914_/X _12441_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _11915_/X sky130_fd_sc_hd__mux2_2
XPHY_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12166_/X _12895_/D _07961_/X vssd1 vssd1 vccd1 vccd1 _12895_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _09957_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11846_/X sky130_fd_sc_hd__mux2_1
XPHY_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _12125_/X _11776_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11777_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10728_ _13253_/Q vssd1 vssd1 vccd1 vccd1 _10730_/A sky130_fd_sc_hd__inv_2
XFILLER_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10659_ _08936_/B _10658_/X _09318_/A vssd1 vssd1 vccd1 vccd1 _10659_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ _12517_/CLK _12329_/D vssd1 vssd1 vccd1 vccd1 _12329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07870_ _13033_/Q _07868_/Y _07869_/Y _12898_/Q vssd1 vssd1 vccd1 vccd1 _07870_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06821_ _12019_/X _12018_/X _06815_/X _06816_/X _06820_/X vssd1 vssd1 vccd1 vccd1
+ _06821_/X sky130_fd_sc_hd__o32a_2
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09540_ _09555_/B vssd1 vssd1 vccd1 vccd1 _09540_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_84_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _13254_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_110_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06752_ _12007_/X _12006_/X _12008_/X _06751_/X vssd1 vssd1 vccd1 vccd1 _06754_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_13_wb_clk_i _12328_/CLK vssd1 vssd1 vccd1 vccd1 _12413_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09471_ _09701_/A vssd1 vssd1 vccd1 vccd1 _09471_/X sky130_fd_sc_hd__buf_2
X_06683_ _06678_/X _06679_/X _06680_/Y _06671_/A _06682_/X vssd1 vssd1 vccd1 vccd1
+ _06683_/X sky130_fd_sc_hd__o221a_1
XFILLER_36_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08422_ _08521_/A vssd1 vssd1 vccd1 vccd1 _08433_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08353_ _12804_/Q _11579_/X _08353_/S vssd1 vssd1 vccd1 vccd1 _12804_/D sky130_fd_sc_hd__mux2_1
XFILLER_196_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07304_ _09226_/A vssd1 vssd1 vccd1 vccd1 _07304_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_177_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08284_ _08284_/A vssd1 vssd1 vccd1 vccd1 _08296_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07235_ _11566_/X _07233_/X _13101_/Q _07234_/X vssd1 vssd1 vccd1 vccd1 _13101_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07166_ _11526_/X _07160_/X _13125_/Q _07161_/X vssd1 vssd1 vccd1 vccd1 _13125_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06117_ _12719_/Q vssd1 vssd1 vccd1 vccd1 _06117_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07097_ _07097_/A _07097_/B _07097_/C _07097_/D vssd1 vssd1 vccd1 vccd1 _07098_/B
+ sky130_fd_sc_hd__or4_1
Xoutput540 _11222_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput551 _11223_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_121_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput562 _11224_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__clkbuf_2
X_06048_ _12707_/Q vssd1 vssd1 vccd1 vccd1 _06048_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput573 _11225_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput584 _12557_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput595 _12567_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_120_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09807_ _09823_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09807_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07999_ _12886_/Q _07996_/X _07997_/X _07998_/X vssd1 vssd1 vccd1 vccd1 _12886_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09738_ _13212_/Q vssd1 vssd1 vccd1 vccd1 _09738_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09669_ _09669_/A vssd1 vssd1 vccd1 vccd1 _09669_/Y sky130_fd_sc_hd__inv_2
XPHY_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11700_ _11699_/X _11396_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12392_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12680_ _12682_/CLK _12680_/D _08758_/X vssd1 vssd1 vccd1 vccd1 _12680_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _10501_/X _12930_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11631_/X sky130_fd_sc_hd__mux2_1
XPHY_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11562_ _12819_/Q _10528_/B _11569_/S vssd1 vssd1 vccd1 vccd1 _11562_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10513_ _12587_/Q _07761_/B _07762_/B vssd1 vssd1 vccd1 vccd1 _10513_/X sky130_fd_sc_hd__a21bo_1
XPHY_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11493_ _10349_/Y _09244_/B _11501_/S vssd1 vssd1 vccd1 vccd1 _11493_/X sky130_fd_sc_hd__mux2_1
XPHY_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13232_ _13237_/CLK _13232_/D _06465_/X vssd1 vssd1 vccd1 vccd1 _13232_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10444_ _10444_/A _10444_/B _10444_/C vssd1 vssd1 vccd1 vccd1 _10455_/D sky130_fd_sc_hd__or3_4
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13163_ _13254_/CLK _13163_/D _07032_/X vssd1 vssd1 vccd1 vccd1 _13163_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10375_ _10375_/A vssd1 vssd1 vccd1 vccd1 _10375_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12114_ _12113_/X _12433_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__mux2_1
X_13094_ _12167_/X _13094_/D _07251_/X vssd1 vssd1 vccd1 vccd1 _13094_/Q sky130_fd_sc_hd__dfrtp_1
X_12045_ _06064_/B _06064_/A _12045_/S vssd1 vssd1 vccd1 vccd1 _12045_/X sky130_fd_sc_hd__mux2_4
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12947_ _12951_/CLK _12947_/D vssd1 vssd1 vccd1 vccd1 _12947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12880_/CLK _12878_/D _08016_/X vssd1 vssd1 vccd1 vccd1 _12878_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11829_ _09920_/X _12854_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11829_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_131_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13268_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_105_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07020_ _11058_/A vssd1 vssd1 vccd1 vccd1 _07020_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08971_ _09067_/A vssd1 vssd1 vccd1 vccd1 _08971_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07922_ _12912_/Q _11501_/X _07932_/S vssd1 vssd1 vccd1 vccd1 _12912_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07853_ _13024_/Q _10357_/A _13037_/Q _10393_/A vssd1 vssd1 vccd1 vccd1 _07858_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06804_ _10737_/A _06804_/B vssd1 vssd1 vccd1 vccd1 _06804_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07784_ _07558_/X _07780_/X _12931_/Q _07781_/X _07775_/X vssd1 vssd1 vccd1 vccd1
+ _12931_/D sky130_fd_sc_hd__a221o_1
XFILLER_65_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06735_ _13205_/Q vssd1 vssd1 vccd1 vccd1 _06735_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09523_ _13174_/Q vssd1 vssd1 vccd1 vccd1 _09524_/A sky130_fd_sc_hd__inv_2
XFILLER_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09454_ _12929_/Q _09438_/X _12925_/Q _09442_/X vssd1 vssd1 vccd1 vccd1 _09454_/X
+ sky130_fd_sc_hd__a22o_1
X_06666_ _12050_/X _12049_/X _06664_/X vssd1 vssd1 vccd1 vccd1 _06666_/X sky130_fd_sc_hd__a21bo_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08405_ _08405_/A vssd1 vssd1 vccd1 vccd1 _08405_/X sky130_fd_sc_hd__clkbuf_1
X_09385_ _12410_/D vssd1 vssd1 vccd1 vccd1 _09385_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06597_ _06602_/A _06602_/B vssd1 vssd1 vccd1 vccd1 _06598_/B sky130_fd_sc_hd__and2_1
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08336_ _08339_/A vssd1 vssd1 vccd1 vccd1 _08336_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08267_ _12836_/Q _08251_/A _07313_/X _08250_/A vssd1 vssd1 vccd1 vccd1 _12836_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07218_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07218_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08198_ _13108_/Q vssd1 vssd1 vccd1 vccd1 _08198_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07149_ _11533_/X _07145_/X _13132_/Q _07146_/X vssd1 vssd1 vccd1 vccd1 _13132_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10160_ _12778_/Q vssd1 vssd1 vccd1 vccd1 _10160_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput370 _11156_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__clkbuf_2
Xoutput381 _11166_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput392 _11176_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10091_ _08273_/Y _10090_/X _08109_/Y _10047_/B vssd1 vssd1 vccd1 vccd1 _10091_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_126_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ _12801_/CLK _12801_/D _08364_/X vssd1 vssd1 vccd1 vccd1 _12801_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_28_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10993_ _12541_/Q _12353_/Q vssd1 vssd1 vccd1 vccd1 _10993_/X sky130_fd_sc_hd__or2_1
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12732_ _12735_/CLK _12732_/D _08621_/X vssd1 vssd1 vccd1 vccd1 _12732_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12664_/CLK _12663_/D _08813_/X vssd1 vssd1 vccd1 vccd1 _12663_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _12968_/Q _12981_/Q _12601_/Q vssd1 vssd1 vccd1 vccd1 _11614_/X sky130_fd_sc_hd__mux2_1
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _12975_/CLK _12594_/D vssd1 vssd1 vccd1 vccd1 _12594_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11545_ _12834_/Q _10793_/B _11546_/S vssd1 vssd1 vccd1 vccd1 _11545_/X sky130_fd_sc_hd__mux2_1
XPHY_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11476_ _12919_/Q _10794_/D _11481_/S vssd1 vssd1 vccd1 vccd1 _11476_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13215_ _13217_/CLK _13215_/D _06629_/X vssd1 vssd1 vccd1 vccd1 _13215_/Q sky130_fd_sc_hd__dfrtp_1
X_10427_ _12813_/Q vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__inv_2
XFILLER_136_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10358_ _10368_/D vssd1 vssd1 vccd1 vccd1 _10360_/B sky130_fd_sc_hd__inv_2
X_13146_ _13146_/CLK _13146_/D _07083_/X vssd1 vssd1 vccd1 vccd1 _13146_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_152_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13077_ _13081_/CLK _13077_/D _07298_/X vssd1 vssd1 vccd1 vccd1 _13077_/Q sky130_fd_sc_hd__dfrtp_4
X_10289_ _10284_/Y _10163_/A _10285_/Y _10165_/A _10288_/X vssd1 vssd1 vccd1 vccd1
+ _10289_/X sky130_fd_sc_hd__o221a_1
X_12028_ _11069_/X _11064_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12028_/X sky130_fd_sc_hd__mux2_2
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06520_ _06520_/A _06520_/B vssd1 vssd1 vccd1 vccd1 _06520_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06451_ _06451_/A vssd1 vssd1 vccd1 vccd1 _06451_/Y sky130_fd_sc_hd__inv_2
X_09170_ _11623_/X _09163_/X _12498_/Q _09164_/X vssd1 vssd1 vccd1 vccd1 _12498_/D
+ sky130_fd_sc_hd__a22o_1
X_06382_ _08504_/A vssd1 vssd1 vccd1 vccd1 _06382_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08121_ _13124_/Q vssd1 vssd1 vccd1 vccd1 _08121_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08052_ _12865_/Q _08040_/X _07296_/X _08041_/X vssd1 vssd1 vccd1 vccd1 _12865_/D
+ sky130_fd_sc_hd__a22o_1
X_07003_ _07012_/A _07012_/B vssd1 vssd1 vccd1 vccd1 _07003_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08954_ _09318_/A _09314_/A _09311_/A _08954_/D vssd1 vssd1 vccd1 vccd1 _10627_/A
+ sky130_fd_sc_hd__or4_4
Xinput109 la_data_in[48] vssd1 vssd1 vccd1 vccd1 input109/X sky130_fd_sc_hd__buf_1
XFILLER_9_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07905_ _07933_/A vssd1 vssd1 vccd1 vccd1 _07917_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08885_ _08963_/A vssd1 vssd1 vccd1 vccd1 _08897_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07836_ _07794_/Y _10397_/A _07833_/Y _12915_/Q _07835_/X vssd1 vssd1 vccd1 vccd1
+ _07836_/X sky130_fd_sc_hd__o221a_1
XFILLER_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07767_ _07769_/A vssd1 vssd1 vccd1 vccd1 _07768_/A sky130_fd_sc_hd__inv_2
XFILLER_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09506_ _09504_/A _09504_/B _09492_/X vssd1 vssd1 vccd1 vccd1 _09506_/Y sky130_fd_sc_hd__o21ai_1
X_06718_ _06750_/A vssd1 vssd1 vccd1 vccd1 _06718_/X sky130_fd_sc_hd__clkbuf_1
X_07698_ _07705_/A vssd1 vssd1 vccd1 vccd1 _07698_/X sky130_fd_sc_hd__buf_2
XFILLER_25_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09437_ _09437_/A vssd1 vssd1 vccd1 vccd1 _09438_/A sky130_fd_sc_hd__inv_2
X_06649_ _06649_/A vssd1 vssd1 vccd1 vccd1 _13215_/D sky130_fd_sc_hd__inv_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09368_ _12415_/Q vssd1 vssd1 vccd1 vccd1 _09368_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08319_ _12819_/Q _11594_/X _08321_/S vssd1 vssd1 vccd1 vccd1 _12819_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09299_ _12942_/Q _10527_/C vssd1 vssd1 vccd1 vccd1 _09299_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11330_ vssd1 vssd1 vccd1 vccd1 _11330_/HI _11330_/LO sky130_fd_sc_hd__conb_1
XFILLER_138_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11261_ vssd1 vssd1 vccd1 vccd1 _11261_/HI _11261_/LO sky130_fd_sc_hd__conb_1
XFILLER_181_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13000_ _13001_/CLK _13000_/D vssd1 vssd1 vccd1 vccd1 _13000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10212_ _10211_/Y _10045_/A _08471_/Y _10113_/A vssd1 vssd1 vccd1 vccd1 _10212_/X
+ sky130_fd_sc_hd__o22a_1
X_11192_ vssd1 vssd1 vccd1 vccd1 _11192_/HI _11192_/LO sky130_fd_sc_hd__conb_1
XFILLER_122_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10143_ _12627_/Q vssd1 vssd1 vccd1 vccd1 _10143_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10074_ _07850_/Y _10070_/X _10073_/X vssd1 vssd1 vccd1 vccd1 _10074_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10976_ _10976_/A _10976_/B vssd1 vssd1 vccd1 vccd1 _10977_/C sky130_fd_sc_hd__or2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12715_ _12717_/CLK _12715_/D _08665_/X vssd1 vssd1 vccd1 vccd1 _12715_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12646_ _12646_/CLK _12646_/D _08856_/X vssd1 vssd1 vccd1 vccd1 _12646_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12577_ _12577_/CLK _12577_/D vssd1 vssd1 vccd1 vccd1 _12577_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _12817_/Q _10528_/C _11533_/S vssd1 vssd1 vccd1 vccd1 _11528_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11459_ _12902_/Q _09243_/D _11459_/S vssd1 vssd1 vccd1 vccd1 _11459_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13129_ _12168_/X _13129_/D _07155_/X vssd1 vssd1 vccd1 vccd1 _13129_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08670_ _08685_/A vssd1 vssd1 vccd1 vccd1 _08670_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07621_ _12947_/Q vssd1 vssd1 vccd1 vccd1 _07678_/A sky130_fd_sc_hd__buf_2
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07552_ _07552_/A vssd1 vssd1 vccd1 vccd1 _07552_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06503_ _13228_/Q vssd1 vssd1 vccd1 vccd1 _06503_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07483_ _07489_/A vssd1 vssd1 vccd1 vccd1 _07483_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09222_ _12469_/Q _09215_/X _07568_/X _09216_/X vssd1 vssd1 vccd1 vccd1 _12469_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06434_ _06886_/A vssd1 vssd1 vccd1 vccd1 _06841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09153_ _09155_/A vssd1 vssd1 vccd1 vccd1 _09163_/A sky130_fd_sc_hd__buf_2
X_06365_ _13252_/Q vssd1 vssd1 vccd1 vccd1 _06365_/X sky130_fd_sc_hd__buf_2
XFILLER_175_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08104_ _12845_/Q _08082_/A _07313_/X _08083_/A vssd1 vssd1 vccd1 vccd1 _12845_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09084_ _12544_/Q _09079_/Y _09180_/D _09083_/X vssd1 vssd1 vccd1 vccd1 _12544_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_148_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06296_ _06269_/X _06281_/X _06295_/Y _13266_/Q _06273_/X vssd1 vssd1 vccd1 vccd1
+ _13266_/D sky130_fd_sc_hd__a32o_1
XFILLER_163_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08035_ _12872_/Q _08024_/X _07990_/X _08026_/X vssd1 vssd1 vccd1 vccd1 _12872_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput80 la_data_in[21] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__buf_1
XFILLER_162_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput91 la_data_in[31] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__buf_1
XFILLER_101_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09986_ _11969_/S _09986_/B _11967_/S _09986_/D vssd1 vssd1 vccd1 vccd1 _10168_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_107_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08937_ _12436_/Q vssd1 vssd1 vccd1 vccd1 _08940_/A sky130_fd_sc_hd__inv_2
XFILLER_112_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08868_ _08963_/A vssd1 vssd1 vccd1 vccd1 _08882_/A sky130_fd_sc_hd__buf_2
XFILLER_57_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07819_ _07819_/A _07819_/B _07819_/C _07818_/X vssd1 vssd1 vccd1 vccd1 _07880_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_45_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08799_ _08798_/X _08781_/X _06271_/Y _12669_/Q _08567_/X vssd1 vssd1 vccd1 vccd1
+ _12669_/D sky130_fd_sc_hd__a32o_1
XFILLER_199_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10830_ _12517_/Q _12329_/Q vssd1 vssd1 vccd1 vccd1 _10830_/X sky130_fd_sc_hd__or2_1
XFILLER_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10761_ _12195_/X vssd1 vssd1 vccd1 vccd1 _10761_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _13243_/CLK _12500_/D vssd1 vssd1 vccd1 vccd1 _12500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10692_ _13240_/Q vssd1 vssd1 vccd1 vccd1 _10693_/A sky130_fd_sc_hd__inv_2
XFILLER_197_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12431_ _12434_/CLK _12431_/D vssd1 vssd1 vccd1 vccd1 _12431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12362_ _12376_/CLK _12362_/D vssd1 vssd1 vccd1 vccd1 _12362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11313_ vssd1 vssd1 vccd1 vccd1 _11313_/HI _11313_/LO sky130_fd_sc_hd__conb_1
XFILLER_5_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12293_ _12296_/CLK _12293_/D vssd1 vssd1 vccd1 vccd1 _12293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11244_ vssd1 vssd1 vccd1 vccd1 _11244_/HI _11244_/LO sky130_fd_sc_hd__conb_1
XFILLER_106_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11175_ vssd1 vssd1 vccd1 vccd1 _11175_/HI _11175_/LO sky130_fd_sc_hd__conb_1
XFILLER_110_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ _10792_/D _10035_/A _08561_/Y _10125_/Y _10140_/A vssd1 vssd1 vccd1 vccd1
+ _10126_/X sky130_fd_sc_hd__o32a_1
XFILLER_121_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10057_ _12878_/Q vssd1 vssd1 vccd1 vccd1 _10057_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10959_ _10958_/A _10958_/B _10958_/Y vssd1 vssd1 vccd1 vccd1 _10977_/B sky130_fd_sc_hd__a21o_1
XFILLER_189_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12629_ _13154_/CLK _12629_/D _08897_/X vssd1 vssd1 vccd1 vccd1 _12629_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_38_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12577_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06150_ _06046_/A _06046_/B _06147_/Y _06149_/Y vssd1 vssd1 vccd1 vccd1 _06151_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_106_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06081_ _12730_/Q _12698_/Q _12730_/Q _12698_/Q vssd1 vssd1 vccd1 vccd1 _06180_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_176_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09840_ _09839_/A _09839_/B _09839_/X vssd1 vssd1 vccd1 vccd1 _09847_/B sky130_fd_sc_hd__a21bo_1
XFILLER_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09771_ _09743_/Y _09745_/Y _09762_/Y vssd1 vssd1 vccd1 vccd1 _09771_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_85_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06983_ _11075_/A _06983_/B vssd1 vssd1 vccd1 vccd1 _06983_/Y sky130_fd_sc_hd__nand2_1
X_08722_ _11827_/X _08715_/X _12693_/Q _08716_/X vssd1 vssd1 vccd1 vccd1 _12693_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ _08653_/A vssd1 vssd1 vccd1 vccd1 _08653_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_93_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07604_ _07611_/A vssd1 vssd1 vccd1 vccd1 _07610_/A sky130_fd_sc_hd__inv_2
XFILLER_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _11956_/X _08575_/X _12747_/Q _08578_/X vssd1 vssd1 vccd1 vccd1 _12747_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07535_ _09019_/B _07531_/X _09185_/A _07532_/X _09023_/A vssd1 vssd1 vccd1 vccd1
+ _13001_/D sky130_fd_sc_hd__o221a_1
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07466_ _11461_/X _07459_/X _13020_/Q _07460_/X vssd1 vssd1 vccd1 vccd1 _13020_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09205_ _12482_/Q _09199_/X _10528_/C _09200_/X vssd1 vssd1 vccd1 vccd1 _12482_/D
+ sky130_fd_sc_hd__a22o_1
X_06417_ _06465_/A vssd1 vssd1 vccd1 vccd1 _06417_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07397_ _11420_/X _07384_/X _13044_/Q _07385_/X vssd1 vssd1 vccd1 vccd1 _13044_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ _12497_/Q _09136_/B vssd1 vssd1 vccd1 vccd1 _09137_/B sky130_fd_sc_hd__or2_1
X_06348_ _06416_/A vssd1 vssd1 vccd1 vccd1 _06370_/A sky130_fd_sc_hd__buf_2
XFILLER_182_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09067_ _09067_/A vssd1 vssd1 vccd1 vccd1 _09067_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06279_ _06269_/X _06247_/X _06278_/Y _13269_/Q _06273_/X vssd1 vssd1 vccd1 vccd1
+ _13269_/D sky130_fd_sc_hd__a32o_1
XFILLER_120_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08018_ _08018_/A vssd1 vssd1 vccd1 vccd1 _08018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09969_ _10034_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _10032_/A sky130_fd_sc_hd__or2_2
XFILLER_131_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12980_ _12984_/CLK _12980_/D vssd1 vssd1 vccd1 vccd1 _12980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11931_ _09519_/X _12792_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11931_/X sky130_fd_sc_hd__mux2_2
XFILLER_150_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11862_ _10108_/Y _12316_/Q _12312_/Q vssd1 vssd1 vccd1 vccd1 _11862_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10813_ _12513_/Q _12325_/Q _10809_/X _10810_/Y vssd1 vssd1 vccd1 vccd1 _10821_/C
+ sky130_fd_sc_hd__o2bb2a_2
XPHY_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _12143_/X _11792_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11793_/X sky130_fd_sc_hd__mux2_1
XPHY_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10744_ _12759_/Q _12758_/Q vssd1 vssd1 vccd1 vccd1 _10744_/Y sky130_fd_sc_hd__nor2_2
XPHY_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10675_ _12437_/Q vssd1 vssd1 vccd1 vccd1 _10675_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12414_ _12995_/CLK _12414_/D vssd1 vssd1 vccd1 vccd1 _12414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12345_ _12570_/CLK _12345_/D vssd1 vssd1 vccd1 vccd1 _12345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12276_ _10231_/X _12902_/Q _11872_/X _10227_/Y _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12292_/D sky130_fd_sc_hd__mux4_2
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11227_ vssd1 vssd1 vccd1 vccd1 _11227_/HI _11227_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11158_ vssd1 vssd1 vccd1 vccd1 _11158_/HI _11158_/LO sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_156_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12570_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10109_ _13077_/Q vssd1 vssd1 vccd1 vccd1 _10109_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11089_ _06368_/X _11045_/A _08535_/A _10742_/X _07030_/X vssd1 vssd1 vccd1 vccd1
+ _11089_/X sky130_fd_sc_hd__a32o_1
XFILLER_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput270 la_oenb[78] vssd1 vssd1 vccd1 vccd1 input270/X sky130_fd_sc_hd__buf_1
Xinput281 la_oenb[88] vssd1 vssd1 vccd1 vccd1 input281/X sky130_fd_sc_hd__buf_1
Xinput292 la_oenb[98] vssd1 vssd1 vccd1 vccd1 input292/X sky130_fd_sc_hd__buf_1
XFILLER_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07320_ _07384_/A vssd1 vssd1 vccd1 vccd1 _07368_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_147_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07251_ _07251_/A vssd1 vssd1 vccd1 vccd1 _07251_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06202_ _06214_/A vssd1 vssd1 vccd1 vccd1 _06202_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_164_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07182_ _11520_/X _07176_/X _13119_/Q _07177_/X vssd1 vssd1 vccd1 vccd1 _13119_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06133_ _06133_/A _06133_/B vssd1 vssd1 vccd1 vccd1 _06134_/A sky130_fd_sc_hd__nand2_1
XFILLER_191_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06064_ _06064_/A _06064_/B vssd1 vssd1 vccd1 vccd1 _06069_/A sky130_fd_sc_hd__nand2_1
XFILLER_172_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09823_ _09823_/A _09823_/B vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__or2_1
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09754_ _09701_/X _09752_/X _09753_/Y _09682_/X vssd1 vssd1 vccd1 vccd1 _09754_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06966_ _06962_/X _06963_/X _06965_/X vssd1 vssd1 vccd1 vccd1 _06966_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08705_ _11834_/X _08700_/X _12700_/Q _08701_/X vssd1 vssd1 vccd1 vccd1 _12700_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09685_ _13238_/Q vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__inv_2
XFILLER_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06897_ _12013_/X vssd1 vssd1 vccd1 vccd1 _06898_/B sky130_fd_sc_hd__inv_2
XFILLER_199_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08636_ _08638_/A vssd1 vssd1 vccd1 vccd1 _08636_/X sky130_fd_sc_hd__clkbuf_1
XPHY_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _08567_/A vssd1 vssd1 vccd1 vccd1 _08567_/X sky130_fd_sc_hd__buf_2
XFILLER_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07518_ _07518_/A vssd1 vssd1 vccd1 vccd1 _07519_/B sky130_fd_sc_hd__buf_2
XPHY_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08498_ _08503_/A vssd1 vssd1 vccd1 vccd1 _08498_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07449_ _11468_/X _07444_/X _13027_/Q _07445_/X vssd1 vssd1 vccd1 vccd1 _13027_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10460_ _10460_/A _10460_/B vssd1 vssd1 vccd1 vccd1 _10462_/A sky130_fd_sc_hd__or2_1
XFILLER_149_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09119_ _12521_/Q _09115_/X _07990_/X _09116_/X vssd1 vssd1 vccd1 vccd1 _12521_/D
+ sky130_fd_sc_hd__a22o_1
X_10391_ _10393_/B vssd1 vssd1 vccd1 vccd1 _10391_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ _12129_/X _12437_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12130_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12061_ _12440_/Q _10678_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _12061_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ _12357_/Q vssd1 vssd1 vccd1 vccd1 _11013_/B sky130_fd_sc_hd__inv_2
XFILLER_2_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12963_ _12975_/CLK _12963_/D vssd1 vssd1 vccd1 vccd1 _12963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11914_ _11913_/X _12441_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11914_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _12166_/X _12894_/D _07964_/X vssd1 vssd1 vccd1 vccd1 _12894_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _09956_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11845_/X sky130_fd_sc_hd__mux2_1
XPHY_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11776_ _09243_/D _11775_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11776_/X sky130_fd_sc_hd__mux2_1
XPHY_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10727_ _13248_/Q _06425_/A _10763_/A _10717_/X _06430_/A vssd1 vssd1 vccd1 vccd1
+ _11145_/A sky130_fd_sc_hd__o221a_1
XFILLER_158_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10658_ _12441_/Q _12442_/Q _12443_/Q vssd1 vssd1 vccd1 vccd1 _10658_/X sky130_fd_sc_hd__o21a_1
XFILLER_167_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10589_ _12403_/D _10594_/A vssd1 vssd1 vccd1 vccd1 _10589_/Y sky130_fd_sc_hd__nor2_1
XFILLER_154_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12328_ _12328_/CLK _12328_/D vssd1 vssd1 vccd1 vccd1 _12328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12259_ _12784_/Q _12857_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12259_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06820_ _06817_/X _06818_/X _12027_/X _06819_/X vssd1 vssd1 vccd1 vccd1 _06820_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_56_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06751_ _12007_/X _12006_/X _12007_/X _12006_/X vssd1 vssd1 vccd1 vccd1 _06751_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06682_ _12199_/X _06688_/B vssd1 vssd1 vccd1 vccd1 _06682_/X sky130_fd_sc_hd__or2_1
X_09470_ _09491_/A vssd1 vssd1 vccd1 vccd1 _09701_/A sky130_fd_sc_hd__buf_2
XFILLER_110_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08421_ _12780_/Q _08417_/X _09242_/A _08418_/X vssd1 vssd1 vccd1 vccd1 _12780_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08352_ _08352_/A vssd1 vssd1 vccd1 vccd1 _08352_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_53_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12999_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07303_ _09185_/C vssd1 vssd1 vccd1 vccd1 _09226_/A sky130_fd_sc_hd__clkbuf_4
X_08283_ _10484_/A _11609_/X _08292_/S vssd1 vssd1 vccd1 vccd1 _12834_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07234_ _07249_/A vssd1 vssd1 vccd1 vccd1 _07234_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07165_ _07167_/A vssd1 vssd1 vccd1 vccd1 _07165_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06116_ _12688_/Q vssd1 vssd1 vccd1 vccd1 _06116_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07096_ _07096_/A _07096_/B _07096_/C _07096_/D vssd1 vssd1 vccd1 vccd1 _07098_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_105_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput530 _11276_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput541 _11286_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__clkbuf_2
X_06047_ _12739_/Q vssd1 vssd1 vccd1 vccd1 _06047_/Y sky130_fd_sc_hd__inv_2
Xoutput552 _11296_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput563 _11306_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__clkbuf_2
XFILLER_121_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput574 _11153_/HI vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__clkbuf_2
Xoutput585 _12558_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput596 _12568_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09806_ _09751_/B _09803_/X _09751_/A _09803_/X _09851_/A vssd1 vssd1 vccd1 vccd1
+ _09808_/B sky130_fd_sc_hd__o221a_1
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07998_ _07998_/A vssd1 vssd1 vccd1 vccd1 _07998_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09737_ _06705_/Y _06710_/Y _09724_/Y _09725_/Y vssd1 vssd1 vccd1 vccd1 _09742_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_27_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06949_ _11077_/A _06954_/B vssd1 vssd1 vccd1 vccd1 _06949_/X sky130_fd_sc_hd__or2_1
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09668_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09669_/A sky130_fd_sc_hd__or2_1
XFILLER_55_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _08623_/A vssd1 vssd1 vccd1 vccd1 _08619_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _13186_/Q _13185_/Q _06905_/Y _06909_/Y vssd1 vssd1 vccd1 vccd1 _09600_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_131_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _10500_/X _12929_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11630_/X sky130_fd_sc_hd__mux2_1
XPHY_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _12818_/Q _09243_/A _11569_/S vssd1 vssd1 vccd1 vccd1 _11561_/X sky130_fd_sc_hd__mux2_1
XPHY_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10512_ _12586_/Q _07760_/B _07761_/B vssd1 vssd1 vccd1 vccd1 _10512_/X sky130_fd_sc_hd__a21bo_1
XFILLER_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11492_ _10345_/X _09243_/C _11492_/S vssd1 vssd1 vccd1 vccd1 _11492_/X sky130_fd_sc_hd__mux2_1
XPHY_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13231_ _13235_/CLK _13231_/D _06478_/X vssd1 vssd1 vccd1 vccd1 _13231_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10443_ _10444_/B _10444_/C _12818_/Q _10442_/B _10437_/X vssd1 vssd1 vccd1 vccd1
+ _10443_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13162_ _13162_/CLK _13162_/D _07034_/X vssd1 vssd1 vccd1 vccd1 _13162_/Q sky130_fd_sc_hd__dfrtp_1
X_10374_ _12913_/Q _10376_/C _10372_/X _10375_/A vssd1 vssd1 vccd1 vccd1 _10374_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12113_ _12433_/Q _12112_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12113_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13093_ _12167_/X _13093_/D _07254_/X vssd1 vssd1 vccd1 vccd1 _13093_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_152_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12044_ _10789_/X _10785_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _12044_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12946_ _12951_/CLK _12946_/D vssd1 vssd1 vccd1 vccd1 _12946_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12877_ _12880_/CLK _12877_/D _08018_/X vssd1 vssd1 vccd1 vccd1 _12877_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11828_ _09918_/Y _12853_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11828_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11759_ _12104_/X _12474_/Q _12103_/S vssd1 vssd1 vccd1 vccd1 _11759_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_100_wb_clk_i _13235_/CLK vssd1 vssd1 vccd1 vccd1 _13223_/CLK sky130_fd_sc_hd__clkbuf_16
X_08970_ _08978_/A vssd1 vssd1 vccd1 vccd1 _09067_/A sky130_fd_sc_hd__buf_6
XFILLER_114_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07921_ _07967_/S vssd1 vssd1 vccd1 vccd1 _07932_/S sky130_fd_sc_hd__buf_2
XFILLER_64_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07852_ _12921_/Q vssd1 vssd1 vccd1 vccd1 _10393_/A sky130_fd_sc_hd__inv_2
XFILLER_84_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06803_ _06806_/A vssd1 vssd1 vccd1 vccd1 _06803_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_110_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07783_ _07536_/X _07780_/X _12932_/Q _07781_/X _07775_/X vssd1 vssd1 vccd1 vccd1
+ _12932_/D sky130_fd_sc_hd__a221o_1
XFILLER_72_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09522_ _09522_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09530_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06734_ _06734_/A _06734_/B vssd1 vssd1 vccd1 vccd1 _06734_/X sky130_fd_sc_hd__or2_1
XFILLER_71_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09453_ _12968_/Q _09440_/X _09450_/X _09452_/X vssd1 vssd1 vccd1 vccd1 _09453_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_80_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06665_ _12048_/X _12047_/X _06664_/X vssd1 vssd1 vccd1 vccd1 _06665_/X sky130_fd_sc_hd__o21a_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08404_ _12787_/Q _08401_/X _07975_/X _08403_/X vssd1 vssd1 vccd1 vccd1 _12787_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09384_ _12405_/D vssd1 vssd1 vccd1 vccd1 _09384_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06596_ _12170_/X _06566_/X _12170_/X _06566_/X vssd1 vssd1 vccd1 vccd1 _06602_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_178_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08335_ _08160_/X _11587_/X _08335_/S vssd1 vssd1 vccd1 vccd1 _12812_/D sky130_fd_sc_hd__mux2_1
XFILLER_193_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08266_ _08282_/A vssd1 vssd1 vccd1 vccd1 _08266_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07217_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07217_/X sky130_fd_sc_hd__clkbuf_1
X_08197_ _13085_/Q vssd1 vssd1 vccd1 vccd1 _08197_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07148_ _07152_/A vssd1 vssd1 vccd1 vccd1 _07148_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07079_ _07069_/X _07074_/X _06346_/Y _13148_/Q _07042_/A vssd1 vssd1 vccd1 vccd1
+ _13148_/D sky130_fd_sc_hd__a32o_1
XFILLER_156_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput371 _11157_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput382 _11167_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10090_ _10090_/A vssd1 vssd1 vccd1 vccd1 _10090_/X sky130_fd_sc_hd__buf_2
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput393 _11177_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12800_ _12890_/CLK _12800_/D _08366_/X vssd1 vssd1 vccd1 vccd1 _12800_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_142_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10992_ _10988_/Y _10991_/X _10988_/Y _10991_/X vssd1 vssd1 vccd1 vccd1 _12352_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_167_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12731_ _12735_/CLK _12731_/D _08623_/X vssd1 vssd1 vccd1 vccd1 _12731_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12664_/CLK _12662_/D _08816_/X vssd1 vssd1 vccd1 vccd1 _12662_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _12967_/Q _12980_/Q _12601_/Q vssd1 vssd1 vccd1 vccd1 _11613_/X sky130_fd_sc_hd__mux2_1
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12593_ _12975_/CLK _12593_/D vssd1 vssd1 vccd1 vccd1 _12593_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ _12833_/Q _10794_/A _11546_/S vssd1 vssd1 vccd1 vccd1 _11544_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11475_ _12918_/Q _10792_/A _11481_/S vssd1 vssd1 vccd1 vccd1 _11475_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13214_ _13217_/CLK _13214_/D _06650_/X vssd1 vssd1 vccd1 vccd1 _13214_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10426_ _08160_/X _10424_/Y _10429_/B _10429_/C _10407_/X vssd1 vssd1 vccd1 vccd1
+ _10426_/X sky130_fd_sc_hd__o221a_1
XFILLER_13_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13145_ _12168_/X _13145_/D _07108_/X vssd1 vssd1 vccd1 vccd1 _13145_/Q sky130_fd_sc_hd__dfrtp_2
X_10357_ _10357_/A _10357_/B _10357_/C vssd1 vssd1 vccd1 vccd1 _10368_/D sky130_fd_sc_hd__or3_4
XFILLER_98_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13076_ _13081_/CLK _13076_/D _07302_/X vssd1 vssd1 vccd1 vccd1 _13076_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10288_ _10286_/Y _10166_/A _10287_/Y _10168_/A vssd1 vssd1 vccd1 vccd1 _10288_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12027_ _11093_/X _11088_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__mux2_4
XFILLER_66_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12929_ _12993_/CLK _12929_/D vssd1 vssd1 vccd1 vccd1 _12929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06450_ _12163_/X vssd1 vssd1 vccd1 vccd1 _06458_/A sky130_fd_sc_hd__inv_2
XFILLER_22_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06381_ _06391_/A vssd1 vssd1 vccd1 vccd1 _06381_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08120_ _12810_/Q vssd1 vssd1 vccd1 vccd1 _10420_/A sky130_fd_sc_hd__inv_2
XFILLER_30_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08051_ _08051_/A vssd1 vssd1 vccd1 vccd1 _08051_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07002_ _06999_/Y _11853_/X _11852_/X _07001_/Y vssd1 vssd1 vccd1 vccd1 _07012_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08953_ _12448_/Q _08953_/B _12140_/S _09316_/A vssd1 vssd1 vccd1 vccd1 _08954_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_9_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07904_ _10388_/A _11508_/X _07904_/S vssd1 vssd1 vccd1 vccd1 _12919_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08884_ _08883_/X _06283_/Y _08878_/X _12635_/Q vssd1 vssd1 vccd1 vccd1 _12635_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07835_ _07814_/Y _07815_/X _13036_/Q _10390_/A vssd1 vssd1 vccd1 vccd1 _07835_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07766_ _12592_/Q _07766_/B vssd1 vssd1 vccd1 vccd1 _07769_/A sky130_fd_sc_hd__or2_1
XFILLER_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ _09521_/A vssd1 vssd1 vccd1 vccd1 _09505_/Y sky130_fd_sc_hd__inv_2
X_06717_ _06658_/X _06710_/Y _06608_/X _06716_/X vssd1 vssd1 vccd1 vccd1 _13207_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07697_ _07688_/Y _07693_/X _07661_/A _07694_/X _07695_/X vssd1 vssd1 vccd1 vccd1
+ _12962_/D sky130_fd_sc_hd__o221a_1
XFILLER_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09436_ _09436_/A vssd1 vssd1 vccd1 vccd1 _09436_/X sky130_fd_sc_hd__clkbuf_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06648_ _06630_/X _06632_/X _06645_/X _06646_/X _06647_/Y vssd1 vssd1 vccd1 vccd1
+ _06649_/A sky130_fd_sc_hd__a32o_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _12406_/Q vssd1 vssd1 vccd1 vccd1 _09367_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06579_ _06579_/A vssd1 vssd1 vccd1 vccd1 _13221_/D sky130_fd_sc_hd__inv_2
XFILLER_123_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08318_ _08325_/A vssd1 vssd1 vccd1 vccd1 _08318_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09298_ _09982_/B vssd1 vssd1 vccd1 vccd1 _10527_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_165_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08249_ _08257_/A vssd1 vssd1 vccd1 vccd1 _08249_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11260_ vssd1 vssd1 vccd1 vccd1 _11260_/HI _11260_/LO sky130_fd_sc_hd__conb_1
XFILLER_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10211_ _12843_/Q vssd1 vssd1 vccd1 vccd1 _10211_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11191_ vssd1 vssd1 vccd1 vccd1 _11191_/HI _11191_/LO sky130_fd_sc_hd__conb_1
XFILLER_137_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10142_ _12882_/Q vssd1 vssd1 vccd1 vccd1 _10142_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10073_ _07885_/Y _10796_/A _08461_/Y _10047_/B vssd1 vssd1 vccd1 vccd1 _10073_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10975_ _11000_/A vssd1 vssd1 vccd1 vccd1 _10975_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12714_ _12717_/CLK _12714_/D _08667_/X vssd1 vssd1 vccd1 vccd1 _12714_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_43_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12645_ _12646_/CLK _12645_/D _08858_/X vssd1 vssd1 vccd1 vccd1 _12645_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12576_ _12576_/CLK _12576_/D vssd1 vssd1 vccd1 vccd1 _12576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11527_ _12816_/Q _09244_/A _11533_/S vssd1 vssd1 vccd1 vccd1 _11527_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11458_ _12901_/Q _09183_/A _11459_/S vssd1 vssd1 vccd1 vccd1 _11458_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10409_ _10405_/Y _08176_/Y _08177_/Y vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__o21a_1
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11389_ _10577_/Y _12400_/D _11392_/S vssd1 vssd1 vccd1 vccd1 _11389_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13128_ _12168_/X _13128_/D _07157_/X vssd1 vssd1 vccd1 vccd1 _13128_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13059_ _12165_/X _13059_/D _07358_/X vssd1 vssd1 vccd1 vccd1 _13059_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07620_ _11611_/X _07610_/A _12966_/Q _07611_/A _07616_/X vssd1 vssd1 vccd1 vccd1
+ _12966_/D sky130_fd_sc_hd__o221a_1
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07551_ _07553_/A vssd1 vssd1 vccd1 vccd1 _07552_/A sky130_fd_sc_hd__inv_2
XFILLER_146_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06502_ _06522_/A vssd1 vssd1 vccd1 vccd1 _06502_/X sky130_fd_sc_hd__clkbuf_1
X_07482_ _11455_/X _07474_/X _13014_/Q _07475_/X vssd1 vssd1 vccd1 vccd1 _13014_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09221_ _12470_/Q _09215_/X _07566_/X _09216_/X vssd1 vssd1 vccd1 vccd1 _12470_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06433_ _06465_/A vssd1 vssd1 vccd1 vccd1 _06433_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ _09152_/A _12307_/D vssd1 vssd1 vccd1 vccd1 _09155_/A sky130_fd_sc_hd__or2_2
X_06364_ _06370_/A vssd1 vssd1 vccd1 vccd1 _06364_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08103_ _08257_/A vssd1 vssd1 vccd1 vccd1 _08103_/X sky130_fd_sc_hd__clkbuf_1
X_09083_ _09083_/A vssd1 vssd1 vccd1 vccd1 _09083_/X sky130_fd_sc_hd__buf_2
X_06295_ _06295_/A vssd1 vssd1 vccd1 vccd1 _06295_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_190_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08034_ _08036_/A vssd1 vssd1 vccd1 vccd1 _08034_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput70 la_data_in[12] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_1
Xinput81 la_data_in[22] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__buf_1
XFILLER_190_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput92 la_data_in[32] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__buf_1
XFILLER_171_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09985_ _12653_/Q vssd1 vssd1 vccd1 vccd1 _09985_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08936_ _08936_/A _08936_/B vssd1 vssd1 vccd1 vccd1 _09318_/A sky130_fd_sc_hd__nand2_2
XFILLER_130_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08867_ _07747_/X _06336_/Y _08837_/A _12641_/Q vssd1 vssd1 vccd1 vccd1 _12641_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07818_ _07799_/Y _07800_/X _13032_/Q _10380_/A _07817_/X vssd1 vssd1 vccd1 vccd1
+ _07818_/X sky130_fd_sc_hd__o221a_1
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08798_ _08814_/A vssd1 vssd1 vccd1 vccd1 _08798_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_8_wb_clk_i _12328_/CLK vssd1 vssd1 vccd1 vccd1 _12852_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07749_ _07749_/A vssd1 vssd1 vccd1 vccd1 _07749_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10760_ _11086_/A vssd1 vssd1 vccd1 vccd1 _10760_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09419_ _12408_/D vssd1 vssd1 vccd1 vccd1 _10599_/B sky130_fd_sc_hd__inv_2
XFILLER_201_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10691_ _10691_/A _10691_/B vssd1 vssd1 vccd1 vccd1 _12185_/S sky130_fd_sc_hd__nor2_8
XFILLER_139_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12430_ _12430_/CLK _12430_/D vssd1 vssd1 vccd1 vccd1 _12430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12361_ _12577_/CLK _12361_/D vssd1 vssd1 vccd1 vccd1 _12361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11312_ vssd1 vssd1 vccd1 vccd1 _11312_/HI _11312_/LO sky130_fd_sc_hd__conb_1
XFILLER_193_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12292_ _12296_/CLK _12292_/D vssd1 vssd1 vccd1 vccd1 _12292_/Q sky130_fd_sc_hd__dfxtp_1
X_11243_ vssd1 vssd1 vccd1 vccd1 _11243_/HI _11243_/LO sky130_fd_sc_hd__conb_1
XFILLER_180_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11174_ vssd1 vssd1 vccd1 vccd1 _11174_/HI _11174_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10125_ _12776_/Q vssd1 vssd1 vccd1 vccd1 _10125_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10056_ _12623_/Q vssd1 vssd1 vccd1 vccd1 _10056_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10958_ _10958_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _10958_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10889_ _12523_/Q _12335_/Q _12522_/Q _12334_/Q vssd1 vssd1 vccd1 vccd1 _10889_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12628_ _13154_/CLK _12628_/D _08901_/X vssd1 vssd1 vccd1 vccd1 _12628_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12559_ _12570_/CLK _12559_/D vssd1 vssd1 vccd1 vccd1 _12559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06080_ _06182_/A _06077_/Y _06079_/Y vssd1 vssd1 vccd1 vccd1 _06133_/A sky130_fd_sc_hd__o21a_1
XFILLER_7_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_78_wb_clk_i _13219_/CLK vssd1 vssd1 vccd1 vccd1 _13213_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09770_ _09770_/A _09803_/A vssd1 vssd1 vccd1 vccd1 _09770_/X sky130_fd_sc_hd__or2_1
X_06982_ _06982_/A vssd1 vssd1 vccd1 vccd1 _11075_/A sky130_fd_sc_hd__buf_2
XFILLER_113_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08721_ _08729_/A vssd1 vssd1 vccd1 vccd1 _08721_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08652_ _11929_/X _08639_/X _12720_/Q _08640_/X vssd1 vssd1 vccd1 vccd1 _12720_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07603_ _12601_/Q _12574_/Q vssd1 vssd1 vccd1 vccd1 _07611_/A sky130_fd_sc_hd__or2_2
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08583_ _08591_/A vssd1 vssd1 vccd1 vccd1 _08583_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07534_ _08978_/A vssd1 vssd1 vccd1 vccd1 _09023_/A sky130_fd_sc_hd__buf_2
XPHY_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07465_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07465_/X sky130_fd_sc_hd__clkbuf_1
X_09204_ _12483_/Q _09199_/X _09243_/A _09200_/X vssd1 vssd1 vccd1 vccd1 _12483_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06416_ _06416_/A vssd1 vssd1 vccd1 vccd1 _06465_/A sky130_fd_sc_hd__clkbuf_2
X_07396_ _07408_/A vssd1 vssd1 vccd1 vccd1 _07396_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09135_ _12496_/Q _09135_/B vssd1 vssd1 vccd1 vccd1 _09136_/B sky130_fd_sc_hd__or2_1
XFILLER_136_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06347_ _07742_/B _06281_/A _06346_/Y _13256_/Q _06306_/A vssd1 vssd1 vccd1 vccd1
+ _13256_/D sky130_fd_sc_hd__a32o_1
XFILLER_194_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09066_ _09067_/A vssd1 vssd1 vccd1 vccd1 _09066_/X sky130_fd_sc_hd__clkbuf_1
X_06278_ _06278_/A vssd1 vssd1 vccd1 vccd1 _06278_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_190_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08017_ _12878_/Q _07996_/A _07309_/X _07998_/A vssd1 vssd1 vccd1 vccd1 _12878_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ _10003_/A vssd1 vssd1 vccd1 vccd1 _09968_/X sky130_fd_sc_hd__buf_4
XFILLER_77_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08919_ _12422_/Q vssd1 vssd1 vccd1 vccd1 _08929_/A sky130_fd_sc_hd__inv_2
XFILLER_170_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09899_ _09896_/Y _09897_/X _06342_/A _09892_/X _09898_/X vssd1 vssd1 vccd1 vccd1
+ _09899_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_100_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11930_ _09509_/Y _12791_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11930_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_0_wb_clk_i clkbuf_opt_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ _10111_/Y _12807_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11861_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _10809_/X _10811_/X _10809_/X _10811_/X vssd1 vssd1 vccd1 vccd1 _12325_/D
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _10528_/C _11791_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11792_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ _10742_/X _10737_/X _06368_/X _10738_/X _10739_/X vssd1 vssd1 vccd1 vccd1
+ _10743_/X sky130_fd_sc_hd__a221o_1
XFILLER_201_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10674_ _08940_/A _08940_/B _09314_/A vssd1 vssd1 vccd1 vccd1 _10674_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_185_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12413_ _12413_/CLK _12413_/D vssd1 vssd1 vccd1 vccd1 _12413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12344_ _12344_/CLK _12344_/D vssd1 vssd1 vccd1 vccd1 _12344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12275_ _10213_/Y _12901_/Q _11871_/X _10207_/Y _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12291_/D sky130_fd_sc_hd__mux4_2
XFILLER_4_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11226_ vssd1 vssd1 vccd1 vccd1 _11226_/HI _11226_/LO sky130_fd_sc_hd__conb_1
XFILLER_49_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11157_ vssd1 vssd1 vccd1 vccd1 _11157_/HI _11157_/LO sky130_fd_sc_hd__conb_1
XFILLER_110_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10108_ _10150_/A _11975_/X vssd1 vssd1 vccd1 vccd1 _10108_/Y sky130_fd_sc_hd__nor2b_1
X_11088_ _10699_/X _11077_/X _06400_/X _11086_/X _11087_/X vssd1 vssd1 vccd1 vccd1
+ _11088_/X sky130_fd_sc_hd__a221o_1
XFILLER_191_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput260 la_oenb[69] vssd1 vssd1 vccd1 vccd1 input260/X sky130_fd_sc_hd__buf_1
Xinput271 la_oenb[79] vssd1 vssd1 vccd1 vccd1 input271/X sky130_fd_sc_hd__buf_1
Xinput282 la_oenb[89] vssd1 vssd1 vccd1 vccd1 input282/X sky130_fd_sc_hd__buf_1
X_10039_ _10792_/D _10151_/A _10036_/Y _10037_/Y _10038_/X vssd1 vssd1 vccd1 vccd1
+ _10039_/X sky130_fd_sc_hd__o32a_1
XFILLER_82_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput293 la_oenb[99] vssd1 vssd1 vccd1 vccd1 input293/X sky130_fd_sc_hd__buf_1
XFILLER_36_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_125_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13279_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07250_ _11560_/X _07248_/X _13095_/Q _07249_/X vssd1 vssd1 vccd1 vccd1 _13095_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06201_ _06195_/Y _06022_/X _06163_/X _06200_/X vssd1 vssd1 vccd1 vccd1 _13283_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_158_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07181_ _07183_/A vssd1 vssd1 vccd1 vccd1 _07181_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06132_ _06182_/A _06132_/B _06132_/C vssd1 vssd1 vccd1 vccd1 _06133_/B sky130_fd_sc_hd__or3_4
XFILLER_184_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06063_ _06063_/A vssd1 vssd1 vccd1 vccd1 _06064_/B sky130_fd_sc_hd__buf_1
XFILLER_144_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09822_ _06503_/Y _09821_/X _06503_/Y _09821_/X vssd1 vssd1 vccd1 vccd1 _09847_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09753_ _09769_/A _09849_/A vssd1 vssd1 vccd1 vccd1 _09753_/Y sky130_fd_sc_hd__nand2_1
X_06965_ _06982_/A _06983_/B vssd1 vssd1 vccd1 vccd1 _06965_/X sky130_fd_sc_hd__or2_1
XFILLER_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08704_ _08714_/A vssd1 vssd1 vccd1 vccd1 _08704_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_95_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09684_ _09684_/A vssd1 vssd1 vccd1 vccd1 _09700_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06896_ _12003_/X _06896_/B vssd1 vssd1 vccd1 vccd1 _06896_/X sky130_fd_sc_hd__or2_1
XFILLER_54_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08635_ _11936_/X _08624_/X _12727_/Q _08625_/X vssd1 vssd1 vccd1 vccd1 _12727_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _08811_/A vssd1 vssd1 vccd1 vccd1 _08567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07517_ _09087_/A vssd1 vssd1 vccd1 vccd1 _07518_/A sky130_fd_sc_hd__inv_2
XFILLER_168_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08497_ _06403_/X _12266_/X _06396_/X _12770_/Q vssd1 vssd1 vccd1 vccd1 _12770_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07448_ _07458_/A vssd1 vssd1 vccd1 vccd1 _07448_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07379_ _07391_/A vssd1 vssd1 vccd1 vccd1 _07379_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09118_ _12522_/Q _09115_/X _07986_/X _09116_/X vssd1 vssd1 vccd1 vccd1 _12522_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10390_ _10390_/A _10390_/B vssd1 vssd1 vccd1 vccd1 _10393_/B sky130_fd_sc_hd__or2_1
XFILLER_198_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09049_ _09051_/A _12156_/X vssd1 vssd1 vccd1 vccd1 _12567_/D sky130_fd_sc_hd__nor2b_1
XFILLER_124_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ _12059_/X _12439_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12060_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11011_ _11013_/A _11010_/A _12356_/Q _11010_/Y vssd1 vssd1 vccd1 vccd1 _12356_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12962_ _12975_/CLK _12962_/D vssd1 vssd1 vccd1 vccd1 _12962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11913_ _12441_/Q _11912_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _11913_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12893_ _12166_/X _12893_/D _07966_/X vssd1 vssd1 vccd1 vccd1 _12893_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11844_ _09955_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11844_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _12125_/X _12478_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11775_/X sky130_fd_sc_hd__mux2_1
XPHY_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10726_ _13248_/Q vssd1 vssd1 vccd1 vccd1 _10763_/A sky130_fd_sc_hd__inv_2
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10657_ _12441_/Q _12442_/Q vssd1 vssd1 vccd1 vccd1 _10657_/X sky130_fd_sc_hd__and2_1
XFILLER_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10588_ _10588_/A vssd1 vssd1 vccd1 vccd1 _11403_/S sky130_fd_sc_hd__inv_2
XFILLER_177_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12327_ _12849_/CLK _12327_/D vssd1 vssd1 vccd1 vccd1 _12327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12258_ _12257_/X _12649_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12258_/X sky130_fd_sc_hd__mux2_2
XFILLER_170_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11209_ vssd1 vssd1 vccd1 vccd1 _11209_/HI _11209_/LO sky130_fd_sc_hd__conb_1
X_12189_ _11110_/A _11051_/A _12199_/S vssd1 vssd1 vccd1 vccd1 _12189_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06750_ _06750_/A vssd1 vssd1 vccd1 vccd1 _06750_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06681_ _06678_/X _06679_/X _06678_/X _06679_/X vssd1 vssd1 vccd1 vccd1 _06688_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_58_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08420_ _08420_/A vssd1 vssd1 vccd1 vccd1 _08420_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08351_ _10405_/A _11580_/X _08353_/S vssd1 vssd1 vccd1 vccd1 _12805_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07302_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07302_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08282_ _08282_/A vssd1 vssd1 vccd1 vccd1 _08282_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07233_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07233_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_93_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _13158_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12474_/CLK sky130_fd_sc_hd__clkbuf_16
X_07164_ _11527_/X _07160_/X _13126_/Q _07161_/X vssd1 vssd1 vccd1 vccd1 _13126_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06115_ _12720_/Q vssd1 vssd1 vccd1 vccd1 _06115_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07095_ _09041_/A _07095_/B vssd1 vssd1 vccd1 vccd1 _07099_/C sky130_fd_sc_hd__or2_1
Xoutput520 _11267_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__clkbuf_2
Xoutput531 _11277_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__clkbuf_2
X_06046_ _06046_/A _06046_/B _06209_/B vssd1 vssd1 vccd1 vccd1 _06197_/B sky130_fd_sc_hd__or3_4
Xoutput542 _11287_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput553 _11297_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__clkbuf_2
Xoutput564 _11307_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput575 _12283_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput586 _12284_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput597 _12285_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09805_ _09771_/Y _09824_/A _09804_/Y vssd1 vssd1 vccd1 vccd1 _09851_/A sky130_fd_sc_hd__o21a_1
XFILLER_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07997_ _09243_/D vssd1 vssd1 vccd1 vccd1 _07997_/X sky130_fd_sc_hd__buf_4
XFILLER_80_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09736_ _09722_/X _09726_/X _09721_/Y _09727_/X vssd1 vssd1 vccd1 vccd1 _09745_/A
+ sky130_fd_sc_hd__o22a_4
X_06948_ _06946_/X _06947_/X _06946_/X _06947_/X vssd1 vssd1 vccd1 vccd1 _06954_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09667_ _13200_/Q _09666_/A _09665_/Y _09666_/Y vssd1 vssd1 vccd1 vccd1 _09668_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06879_ _06879_/A vssd1 vssd1 vccd1 vccd1 _06883_/A sky130_fd_sc_hd__inv_2
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _11943_/X _08608_/X _12734_/Q _08610_/X vssd1 vssd1 vccd1 vccd1 _12734_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _12872_/Q vssd1 vssd1 vccd1 vccd1 _09598_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08569_/A vssd1 vssd1 vccd1 vccd1 _08549_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ _12817_/Q _10528_/C _11569_/S vssd1 vssd1 vccd1 vccd1 _11560_/X sky130_fd_sc_hd__mux2_1
XFILLER_196_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10511_ _12585_/Q _07759_/B _07760_/B vssd1 vssd1 vccd1 vccd1 _10511_/X sky130_fd_sc_hd__a21bo_1
XPHY_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11491_ _10344_/Y _09243_/D _11492_/S vssd1 vssd1 vccd1 vccd1 _11491_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13236_/CLK _13230_/D _06482_/X vssd1 vssd1 vccd1 vccd1 _13230_/Q sky130_fd_sc_hd__dfrtp_1
X_10442_ _10458_/A _10442_/B _10442_/C vssd1 vssd1 vccd1 vccd1 _10442_/Y sky130_fd_sc_hd__nor3_1
XFILLER_148_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13161_ _13161_/CLK _13161_/D _07044_/X vssd1 vssd1 vccd1 vccd1 _13161_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_164_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10373_ _10373_/A _10373_/B vssd1 vssd1 vccd1 vccd1 _10375_/A sky130_fd_sc_hd__or2_1
XFILLER_163_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12112_ _10670_/Y _12433_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12112_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13092_ _12167_/X _13092_/D _07256_/X vssd1 vssd1 vccd1 vccd1 _13092_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12043_ _10787_/Y _10783_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _12043_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12945_ _13241_/CLK _12945_/D _07728_/X vssd1 vssd1 vccd1 vccd1 _12945_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12876_ _12892_/CLK _12876_/D _08021_/X vssd1 vssd1 vccd1 vccd1 _12876_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _09913_/X _12852_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11827_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11757_/X _12100_/X _11774_/S vssd1 vssd1 vccd1 vccd1 _12429_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10709_ _13239_/Q _11107_/A _10686_/A _11100_/A _06470_/Y vssd1 vssd1 vccd1 vccd1
+ _11079_/A sky130_fd_sc_hd__o221a_1
XPHY_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11689_ _11398_/X _09243_/A _11691_/S vssd1 vssd1 vccd1 vccd1 _11689_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07920_ _07931_/A vssd1 vssd1 vccd1 vccd1 _07920_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07851_ _13032_/Q _10380_/A _07850_/Y _12894_/Q vssd1 vssd1 vccd1 vccd1 _07858_/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_140_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12880_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_96_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06802_ _06658_/X _06796_/Y _06769_/X _06801_/X vssd1 vssd1 vccd1 vccd1 _13198_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_84_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_1
X_07782_ _07545_/X _07780_/X _12933_/Q _07781_/X _07775_/X vssd1 vssd1 vccd1 vccd1
+ _12933_/D sky130_fd_sc_hd__a221o_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09521_ _09521_/A _09521_/B vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__or2_1
X_06733_ _11989_/X _06702_/X _11989_/X _06702_/X vssd1 vssd1 vccd1 vccd1 _06734_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09452_ _12980_/Q _09436_/X _12996_/Q _09451_/X vssd1 vssd1 vccd1 vccd1 _09452_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06664_ _12050_/X _12049_/X vssd1 vssd1 vccd1 vccd1 _06664_/X sky130_fd_sc_hd__or2_1
XFILLER_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _08418_/A vssd1 vssd1 vccd1 vccd1 _08403_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09383_ _12407_/D vssd1 vssd1 vccd1 vccd1 _10599_/A sky130_fd_sc_hd__inv_2
X_06595_ _06588_/X _06592_/X _06598_/A vssd1 vssd1 vccd1 vccd1 _06602_/A sky130_fd_sc_hd__a21oi_2
X_08334_ _08339_/A vssd1 vssd1 vccd1 vccd1 _08334_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08265_ _12837_/Q _08251_/A _07309_/X _08250_/A vssd1 vssd1 vccd1 vccd1 _12837_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07216_ _11573_/X _07201_/X _13108_/Q _07204_/X vssd1 vssd1 vccd1 vccd1 _13108_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08196_ _08193_/Y _12834_/Q _08194_/Y _12806_/Q _08195_/X vssd1 vssd1 vccd1 vccd1
+ _08209_/A sky130_fd_sc_hd__a221o_1
XFILLER_118_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07147_ _11534_/X _07145_/X _13133_/Q _07146_/X vssd1 vssd1 vccd1 vccd1 _13133_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07078_ _07078_/A vssd1 vssd1 vccd1 vccd1 _07078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput372 _11158_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__clkbuf_2
X_06029_ _12746_/Q _12714_/Q _12746_/Q _12714_/Q vssd1 vssd1 vccd1 vccd1 _06029_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_121_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput383 _11168_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__clkbuf_2
Xoutput394 _11178_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09719_ _09747_/A _09825_/A vssd1 vssd1 vccd1 vccd1 _09719_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10991_ _10975_/Y _10983_/Y _10980_/Y _10990_/X vssd1 vssd1 vccd1 vccd1 _10991_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_56_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12730_ _12735_/CLK _12730_/D _08628_/X vssd1 vssd1 vccd1 vccd1 _12730_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12661_ _12664_/CLK _12661_/D _08819_/X vssd1 vssd1 vccd1 vccd1 _12661_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _12966_/Q _12979_/Q _12601_/Q vssd1 vssd1 vccd1 vccd1 _11612_/X sky130_fd_sc_hd__mux2_1
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12937_/CLK _12592_/D vssd1 vssd1 vccd1 vccd1 _12592_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ _12832_/Q _10794_/B _11543_/S vssd1 vssd1 vccd1 vccd1 _11543_/X sky130_fd_sc_hd__mux2_1
XPHY_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11474_ _12917_/Q _10792_/B _11481_/S vssd1 vssd1 vccd1 vccd1 _11474_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13213_ _13213_/CLK _13213_/D _06657_/X vssd1 vssd1 vccd1 vccd1 _13213_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10425_ _12812_/Q vssd1 vssd1 vccd1 vccd1 _10429_/B sky130_fd_sc_hd__inv_2
XFILLER_104_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13144_ _12168_/X _13144_/D _07118_/X vssd1 vssd1 vccd1 vccd1 _13144_/Q sky130_fd_sc_hd__dfrtp_1
X_10356_ _10357_/B _10357_/C _12907_/Q _10355_/B _10350_/X vssd1 vssd1 vccd1 vccd1
+ _10356_/X sky130_fd_sc_hd__o221a_1
XFILLER_97_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13075_ _12169_/A0 _13075_/D _07307_/X vssd1 vssd1 vccd1 vccd1 _13075_/Q sky130_fd_sc_hd__dfrtp_1
X_10287_ _12651_/Q vssd1 vssd1 vccd1 vccd1 _10287_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12026_ _11120_/X _11113_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _12026_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12928_ _12993_/CLK _12928_/D vssd1 vssd1 vccd1 vccd1 _12928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _12890_/CLK _12859_/D _08070_/X vssd1 vssd1 vccd1 vccd1 _12859_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06380_ _06361_/X _12222_/X _06375_/X _06379_/X vssd1 vssd1 vccd1 vccd1 _13248_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08050_ _12866_/Q _08040_/X _07293_/X _08041_/X vssd1 vssd1 vccd1 vccd1 _12866_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07001_ _11853_/X vssd1 vssd1 vccd1 vccd1 _07001_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08952_ _09315_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__or2_2
XFILLER_9_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07903_ _07903_/A vssd1 vssd1 vccd1 vccd1 _07903_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08883_ _08898_/A vssd1 vssd1 vccd1 vccd1 _08883_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07834_ _12920_/Q vssd1 vssd1 vccd1 vccd1 _10390_/A sky130_fd_sc_hd__inv_2
XFILLER_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07765_ _12591_/Q _07765_/B vssd1 vssd1 vccd1 vccd1 _07766_/B sky130_fd_sc_hd__or2_1
XFILLER_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06716_ _06711_/X _06712_/X _06704_/X _06694_/X _06715_/X vssd1 vssd1 vccd1 vccd1
+ _06716_/X sky130_fd_sc_hd__o221a_1
X_09504_ _09504_/A _09504_/B vssd1 vssd1 vccd1 vccd1 _09521_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07696_ _07688_/Y _07693_/X _12963_/Q _07694_/X _07695_/X vssd1 vssd1 vccd1 vccd1
+ _12963_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09435_ _10527_/A _09435_/B _10527_/C vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__and3_1
X_06647_ _13215_/Q vssd1 vssd1 vccd1 vccd1 _06647_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09366_ _12463_/Q vssd1 vssd1 vccd1 vccd1 _09366_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06578_ _06526_/X _06573_/B _06576_/Y _06556_/X _06577_/Y vssd1 vssd1 vccd1 vccd1
+ _06579_/A sky130_fd_sc_hd__o32a_1
XFILLER_200_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08317_ _12820_/Q _11595_/X _08321_/S vssd1 vssd1 vccd1 vccd1 _12820_/D sky130_fd_sc_hd__mux2_1
X_09297_ _12941_/Q vssd1 vssd1 vccd1 vccd1 _09297_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08248_ _12844_/Q _08191_/X _09019_/A _08275_/A vssd1 vssd1 vccd1 vccd1 _12844_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08179_ _08159_/Y _08160_/X _13114_/Q _08176_/Y _08178_/X vssd1 vssd1 vccd1 vccd1
+ _08179_/X sky130_fd_sc_hd__a221o_1
XFILLER_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10210_ _08210_/Y _10151_/X _10209_/X vssd1 vssd1 vccd1 vccd1 _10210_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11190_ vssd1 vssd1 vccd1 vccd1 _11190_/HI _11190_/LO sky130_fd_sc_hd__conb_1
XFILLER_122_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10141_ _10141_/A vssd1 vssd1 vccd1 vccd1 _10141_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10072_ _08226_/Y _10070_/X _10071_/X vssd1 vssd1 vccd1 vccd1 _10072_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10974_ _12538_/Q _12350_/Q _12538_/Q _12350_/Q vssd1 vssd1 vccd1 vccd1 _11000_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12713_ _12713_/CLK _12713_/D _08669_/X vssd1 vssd1 vccd1 vccd1 _12713_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12644_ _12646_/CLK _12644_/D _08860_/X vssd1 vssd1 vccd1 vccd1 _12644_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ _12576_/CLK _12575_/D vssd1 vssd1 vccd1 vccd1 _12575_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11526_ _12815_/Q _09244_/B _11533_/S vssd1 vssd1 vccd1 vccd1 _11526_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11457_ _12900_/Q input358/X _11459_/S vssd1 vssd1 vccd1 vccd1 _11457_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10408_ _10405_/A _12804_/Q _10405_/Y _08176_/Y _10407_/X vssd1 vssd1 vccd1 vccd1
+ _10408_/X sky130_fd_sc_hd__o221a_1
X_11388_ _10580_/X _12401_/D _11390_/S vssd1 vssd1 vccd1 vccd1 _11388_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10339_ _07821_/X _10337_/Y _10342_/B _10342_/C _10320_/X vssd1 vssd1 vccd1 vccd1
+ _10339_/X sky130_fd_sc_hd__o221a_1
X_13127_ _12168_/X _13127_/D _07159_/X vssd1 vssd1 vccd1 vccd1 _13127_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13058_ _12165_/X _13058_/D _07360_/X vssd1 vssd1 vccd1 vccd1 _13058_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12009_ _11117_/X _11105_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _12009_/X sky130_fd_sc_hd__mux2_2
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07550_ _11982_/S _11356_/S vssd1 vssd1 vccd1 vccd1 _07553_/A sky130_fd_sc_hd__nand2_2
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06501_ _06440_/X _06488_/Y _06489_/X _06500_/Y vssd1 vssd1 vccd1 vccd1 _13229_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07481_ _07489_/A vssd1 vssd1 vccd1 vccd1 _07481_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09220_ _12471_/Q _09215_/X _07564_/X _09216_/X vssd1 vssd1 vccd1 vccd1 _12471_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06432_ _06420_/X _06431_/X _06420_/X _13237_/Q vssd1 vssd1 vccd1 vccd1 _13237_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ _12509_/Q _09147_/X _07947_/A _13001_/Q _09150_/X vssd1 vssd1 vccd1 vccd1
+ _11634_/S sky130_fd_sc_hd__o2111ai_4
X_06363_ _06361_/X _12232_/X _06358_/X _06362_/X vssd1 vssd1 vccd1 vccd1 _13253_/D
+ sky130_fd_sc_hd__o22a_1
X_08102_ _12846_/Q _08082_/A _07309_/X _08083_/A vssd1 vssd1 vccd1 vccd1 _12846_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09082_ _12545_/Q _09079_/A _09180_/C _09079_/Y vssd1 vssd1 vccd1 vccd1 _12545_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06294_ _06132_/C _06180_/B _06132_/C _06180_/B vssd1 vssd1 vccd1 vccd1 _06295_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_08033_ _12873_/Q _08024_/X _07986_/X _08026_/X vssd1 vssd1 vccd1 vccd1 _12873_/D
+ sky130_fd_sc_hd__a22o_1
Xinput60 la_data_in[119] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_1
Xinput71 la_data_in[13] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_1
Xinput82 la_data_in[23] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__buf_1
Xinput93 la_data_in[33] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__buf_1
XFILLER_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09984_ _09984_/A _09984_/B _11967_/S _09986_/D vssd1 vssd1 vccd1 vccd1 _10165_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_103_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08935_ _12443_/Q _11916_/S vssd1 vssd1 vccd1 vccd1 _08936_/B sky130_fd_sc_hd__and2b_1
XFILLER_130_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08866_ _08866_/A vssd1 vssd1 vccd1 vccd1 _08866_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater650 _07990_/A vssd1 vssd1 vccd1 vccd1 _09244_/B sky130_fd_sc_hd__buf_8
X_07817_ _07814_/Y _07815_/X _07816_/Y _12902_/Q vssd1 vssd1 vccd1 vccd1 _07817_/X
+ sky130_fd_sc_hd__o22a_1
X_08797_ _12610_/Q vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__clkbuf_2
X_07748_ _12942_/Q _07747_/X _11983_/X vssd1 vssd1 vccd1 vccd1 _12942_/D sky130_fd_sc_hd__mux2_1
XFILLER_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07679_ _07679_/A _07685_/A vssd1 vssd1 vccd1 vccd1 _07680_/A sky130_fd_sc_hd__or2_1
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09418_ _09418_/A vssd1 vssd1 vccd1 vccd1 _10525_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10690_ _11045_/A vssd1 vssd1 vccd1 vccd1 _10691_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_179_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09349_ _12544_/Q vssd1 vssd1 vccd1 vccd1 _09349_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12360_ _13257_/CLK _12360_/D vssd1 vssd1 vccd1 vccd1 _12360_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_139_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11311_ vssd1 vssd1 vccd1 vccd1 _11311_/HI _11311_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12291_ _12296_/CLK _12291_/D vssd1 vssd1 vccd1 vccd1 _12291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11242_ vssd1 vssd1 vccd1 vccd1 _11242_/HI _11242_/LO sky130_fd_sc_hd__conb_1
XFILLER_10_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11173_ vssd1 vssd1 vccd1 vccd1 _11173_/HI _11173_/LO sky130_fd_sc_hd__conb_1
XFILLER_180_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10124_ _12865_/Q vssd1 vssd1 vccd1 vccd1 _10124_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10055_ _13009_/Q _10049_/X _13042_/Q _10051_/X _10054_/Y vssd1 vssd1 vccd1 vccd1
+ _10055_/X sky130_fd_sc_hd__a221o_1
XFILLER_180_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10957_ _12347_/Q vssd1 vssd1 vccd1 vccd1 _10958_/B sky130_fd_sc_hd__inv_2
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10888_ _10890_/A _10890_/B _10888_/C _10888_/D vssd1 vssd1 vccd1 vccd1 _10888_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_148_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ _12765_/CLK _12627_/D _08903_/X vssd1 vssd1 vccd1 vccd1 _12627_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12558_ _12558_/CLK _12558_/D vssd1 vssd1 vccd1 vccd1 _12558_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11509_ _10392_/Y _10794_/C _11513_/S vssd1 vssd1 vccd1 vccd1 _11509_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12489_ _12489_/CLK _12489_/D vssd1 vssd1 vccd1 vccd1 _12489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06981_ _07006_/A vssd1 vssd1 vccd1 vccd1 _06981_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08720_ _11828_/X _08715_/X _12694_/Q _08716_/X vssd1 vssd1 vccd1 vccd1 _12694_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_47_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12455_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_100_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08651_ _08653_/A vssd1 vssd1 vccd1 vccd1 _08651_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07602_ _07609_/A _07602_/B vssd1 vssd1 vccd1 vccd1 _12976_/D sky130_fd_sc_hd__nor2_1
XFILLER_93_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08582_ _11957_/X _08575_/X _12748_/Q _08578_/X vssd1 vssd1 vccd1 vccd1 _12748_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07533_ _08854_/A vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__buf_2
XFILLER_23_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07464_ _11462_/X _07459_/X _13021_/Q _07460_/X vssd1 vssd1 vccd1 vccd1 _13021_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09203_ _12484_/Q _09199_/X _10528_/B _09200_/X vssd1 vssd1 vccd1 vccd1 _12484_/D
+ sky130_fd_sc_hd__a22o_1
X_06415_ _13238_/Q _06415_/B vssd1 vssd1 vccd1 vccd1 _13238_/D sky130_fd_sc_hd__or2_1
XFILLER_148_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07395_ _11421_/X _07384_/X _13045_/Q _07385_/X vssd1 vssd1 vccd1 vccd1 _13045_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09134_ _12495_/Q _12494_/Q vssd1 vssd1 vccd1 vccd1 _09135_/B sky130_fd_sc_hd__or2_1
X_06346_ _06346_/A vssd1 vssd1 vccd1 vccd1 _06346_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_136_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09065_ _09067_/A vssd1 vssd1 vccd1 vccd1 _09065_/X sky130_fd_sc_hd__clkbuf_1
X_06277_ _06075_/A _06276_/X _06075_/A _06276_/X vssd1 vssd1 vccd1 vccd1 _06278_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_68_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08016_ _08018_/A vssd1 vssd1 vccd1 vccd1 _08016_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09967_ _10010_/A vssd1 vssd1 vccd1 vccd1 _10003_/A sky130_fd_sc_hd__buf_2
X_08918_ _12423_/Q vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__inv_2
XFILLER_131_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09898_ _12879_/Q _09910_/B vssd1 vssd1 vccd1 vccd1 _09898_/X sky130_fd_sc_hd__or2_1
XFILLER_85_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08849_ _08849_/A vssd1 vssd1 vccd1 vccd1 _08849_/X sky130_fd_sc_hd__buf_2
XFILLER_73_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11860_ _10089_/Y _12315_/Q _12312_/Q vssd1 vssd1 vccd1 vccd1 _11860_/X sky130_fd_sc_hd__mux2_2
XFILLER_73_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _12513_/Q _12325_/Q _10810_/Y vssd1 vssd1 vccd1 vccd1 _10811_/X sky130_fd_sc_hd__a21o_1
X_11791_ _12143_/X _12482_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11791_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10742_ _10742_/A vssd1 vssd1 vccd1 vccd1 _10742_/X sky130_fd_sc_hd__buf_2
XFILLER_129_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10673_ _08940_/B _10672_/X _09314_/A vssd1 vssd1 vccd1 vccd1 _10673_/X sky130_fd_sc_hd__o21a_1
XFILLER_159_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12412_ _13001_/CLK _12412_/D vssd1 vssd1 vccd1 vccd1 _12412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12343_ _12537_/CLK _12343_/D vssd1 vssd1 vccd1 vccd1 _12343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12274_ _10194_/Y _12900_/Q _11869_/X _11870_/X _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12290_/D sky130_fd_sc_hd__mux4_2
XFILLER_141_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11225_ vssd1 vssd1 vccd1 vccd1 _11225_/HI _11225_/LO sky130_fd_sc_hd__conb_1
XFILLER_150_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11156_ vssd1 vssd1 vccd1 vccd1 _11156_/HI _11156_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10107_ _10107_/A _10107_/B _10107_/C _10107_/D vssd1 vssd1 vccd1 vccd1 _10107_/Y
+ sky130_fd_sc_hd__nand4_2
X_11087_ _12195_/X vssd1 vssd1 vccd1 vccd1 _11087_/X sky130_fd_sc_hd__clkbuf_2
Xinput250 la_oenb[5] vssd1 vssd1 vccd1 vccd1 input250/X sky130_fd_sc_hd__buf_1
Xinput261 la_oenb[6] vssd1 vssd1 vccd1 vccd1 input261/X sky130_fd_sc_hd__buf_1
Xinput272 la_oenb[7] vssd1 vssd1 vccd1 vccd1 input272/X sky130_fd_sc_hd__buf_1
X_10038_ _10140_/A vssd1 vssd1 vccd1 vccd1 _10038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput283 la_oenb[8] vssd1 vssd1 vccd1 vccd1 input283/X sky130_fd_sc_hd__buf_1
Xinput294 la_oenb[9] vssd1 vssd1 vccd1 vccd1 input294/X sky130_fd_sc_hd__buf_1
XFILLER_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11989_ _11125_/X _11118_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _11989_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_165_wb_clk_i clkbuf_opt_1_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12296_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06200_ _06029_/Y _06199_/Y _06029_/Y _06199_/Y vssd1 vssd1 vccd1 vccd1 _06200_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_13_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07180_ _11521_/X _07176_/X _13120_/Q _07177_/X vssd1 vssd1 vccd1 vccd1 _13120_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06131_ _06130_/A _06094_/X _06096_/X _06130_/X vssd1 vssd1 vccd1 vccd1 _06132_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_117_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06062_ _12733_/Q _12701_/Q vssd1 vssd1 vccd1 vccd1 _06063_/A sky130_fd_sc_hd__or2_1
XFILLER_105_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09821_ _06508_/Y _09820_/X _06508_/Y _09820_/X vssd1 vssd1 vccd1 vccd1 _09821_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09752_ _09769_/A _09849_/A vssd1 vssd1 vccd1 vccd1 _09752_/X sky130_fd_sc_hd__or2_1
XFILLER_100_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06964_ _06962_/X _06963_/X _06962_/X _06963_/X vssd1 vssd1 vccd1 vccd1 _06983_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08703_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08714_/A sky130_fd_sc_hd__clkbuf_2
X_09683_ _09471_/X _09677_/X _09678_/Y _09682_/X vssd1 vssd1 vccd1 vccd1 _09683_/X
+ sky130_fd_sc_hd__a31o_1
X_06895_ _12000_/X _06876_/X _12000_/X _06876_/X vssd1 vssd1 vccd1 vccd1 _06896_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08634_ _08638_/A vssd1 vssd1 vccd1 vccd1 _08634_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08781_/A vssd1 vssd1 vccd1 vccd1 _08565_/X sky130_fd_sc_hd__buf_2
XPHY_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07516_ _10527_/A _10527_/B _09986_/B vssd1 vssd1 vccd1 vccd1 _09087_/A sky130_fd_sc_hd__or3_4
XPHY_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08496_ _08503_/A vssd1 vssd1 vccd1 vccd1 _08496_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07447_ _07462_/A vssd1 vssd1 vccd1 vccd1 _07458_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07378_ _07462_/A vssd1 vssd1 vccd1 vccd1 _07391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09117_ _12523_/Q _09115_/X _07983_/X _09116_/X vssd1 vssd1 vccd1 vccd1 _12523_/D
+ sky130_fd_sc_hd__a22o_1
X_06329_ _06344_/A vssd1 vssd1 vccd1 vccd1 _06329_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ _09051_/A _12157_/X vssd1 vssd1 vccd1 vccd1 _12568_/D sky130_fd_sc_hd__nor2b_1
XFILLER_190_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11010_ _11010_/A vssd1 vssd1 vccd1 vccd1 _11010_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12961_ _12961_/CLK _12961_/D vssd1 vssd1 vccd1 vccd1 _12961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11912_ _11911_/X _12441_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _11912_/X sky130_fd_sc_hd__mux2_1
XPHY_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _12892_/CLK _12892_/D _07968_/X vssd1 vssd1 vccd1 vccd1 _12892_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _09954_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11843_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11774_ _11773_/X _12115_/X _11774_/S vssd1 vssd1 vccd1 vccd1 _12433_/D sky130_fd_sc_hd__mux2_1
XPHY_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10725_ _13249_/Q _06425_/A _10758_/A _10717_/X _06430_/X vssd1 vssd1 vccd1 vccd1
+ _10790_/A sky130_fd_sc_hd__o221a_1
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10656_ _12441_/Q vssd1 vssd1 vccd1 vccd1 _10656_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10587_ _12403_/D _12406_/D _10586_/B _10594_/A vssd1 vssd1 vccd1 vccd1 _10588_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_166_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12326_ _12999_/CLK _12326_/D vssd1 vssd1 vccd1 vccd1 _12326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12257_ _12783_/Q _12856_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12257_/X sky130_fd_sc_hd__mux2_1
X_11208_ vssd1 vssd1 vccd1 vccd1 _11208_/HI _11208_/LO sky130_fd_sc_hd__conb_1
XFILLER_123_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12188_ _10708_/X _11079_/A _12202_/S vssd1 vssd1 vccd1 vccd1 _12188_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11139_ _11139_/A vssd1 vssd1 vccd1 vccd1 _11139_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06680_ _06680_/A vssd1 vssd1 vccd1 vccd1 _06680_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08350_ _08352_/A vssd1 vssd1 vccd1 vccd1 _08350_/X sky130_fd_sc_hd__clkbuf_1
X_07301_ _13077_/Q _07285_/X _07300_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _13077_/D
+ sky130_fd_sc_hd__a22o_1
X_08281_ _12835_/Q _11610_/X _08292_/S vssd1 vssd1 vccd1 vccd1 _12835_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07232_ _07236_/A vssd1 vssd1 vccd1 vccd1 _07232_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07163_ _07167_/A vssd1 vssd1 vccd1 vccd1 _07163_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06114_ _12721_/Q _12689_/Q _06112_/Y _06113_/Y vssd1 vssd1 vccd1 vccd1 _06125_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07094_ _07094_/A vssd1 vssd1 vccd1 vccd1 _09071_/B sky130_fd_sc_hd__inv_2
XFILLER_145_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput510 _11258_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput521 _11268_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06045_ _06045_/A _06044_/Y vssd1 vssd1 vccd1 vccd1 _06209_/B sky130_fd_sc_hd__or2b_2
Xoutput532 _11278_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_62_wb_clk_i _12960_/CLK vssd1 vssd1 vccd1 vccd1 _13244_/CLK sky130_fd_sc_hd__clkbuf_16
Xoutput543 _11288_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__clkbuf_2
Xoutput554 _11298_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__clkbuf_2
Xoutput565 _11308_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__clkbuf_2
Xoutput576 _12293_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput587 _12559_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__clkbuf_2
Xoutput598 _12569_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09804_ _09780_/Y _09782_/Y _09790_/Y vssd1 vssd1 vccd1 vccd1 _09804_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07996_ _07996_/A vssd1 vssd1 vccd1 vccd1 _07996_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09735_ _09886_/A _09735_/B vssd1 vssd1 vccd1 vccd1 _09735_/X sky130_fd_sc_hd__or2_1
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06947_ _12005_/X _06928_/X _12005_/X _06928_/X vssd1 vssd1 vccd1 vccd1 _06947_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09666_ _09666_/A vssd1 vssd1 vccd1 vccd1 _09666_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06878_ _11997_/X _11994_/X _06872_/X _06873_/X _06877_/X vssd1 vssd1 vccd1 vccd1
+ _06879_/A sky130_fd_sc_hd__o32a_1
XFILLER_54_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08617_ _08623_/A vssd1 vssd1 vccd1 vccd1 _08617_/X sky130_fd_sc_hd__clkbuf_1
XPHY_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09597_ _09471_/X _09593_/X _09594_/Y _09596_/X vssd1 vssd1 vccd1 vccd1 _09597_/X
+ sky130_fd_sc_hd__a31o_1
XPHY_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08548_/A vssd1 vssd1 vccd1 vccd1 _12752_/D sky130_fd_sc_hd__inv_2
XPHY_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08479_ _13058_/Q _10362_/B _13061_/Q _10367_/A _08478_/X vssd1 vssd1 vccd1 vccd1
+ _08482_/C sky130_fd_sc_hd__o221a_1
XPHY_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10510_ _12584_/Q _07758_/B _07759_/B vssd1 vssd1 vccd1 vccd1 _10510_/X sky130_fd_sc_hd__a21bo_1
XFILLER_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11490_ _10339_/X _09183_/A _11492_/S vssd1 vssd1 vccd1 vccd1 _11490_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10441_ _08187_/X _10439_/C _10439_/A vssd1 vssd1 vccd1 vccd1 _10442_/C sky130_fd_sc_hd__o21a_1
XFILLER_109_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10372_ _10372_/A vssd1 vssd1 vccd1 vccd1 _10372_/X sky130_fd_sc_hd__clkbuf_2
X_13160_ _13161_/CLK _13160_/D _07046_/X vssd1 vssd1 vccd1 vccd1 _13160_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12111_ _12110_/X _12432_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12111_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13091_ _12167_/X _13091_/D _07258_/X vssd1 vssd1 vccd1 vccd1 _13091_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_156_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12042_ _10785_/X _10786_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _12042_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12944_ _13161_/CLK _12944_/D _07734_/X vssd1 vssd1 vccd1 vccd1 _12944_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _12875_/CLK _12875_/D _08028_/X vssd1 vssd1 vccd1 vccd1 _12875_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _09911_/Y _12851_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11826_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11757_ _12100_/X _11756_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11757_/X sky130_fd_sc_hd__mux2_1
XPHY_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10708_ _06407_/X _11107_/A _10693_/X _11100_/A _06470_/Y vssd1 vssd1 vccd1 vccd1
+ _10708_/X sky130_fd_sc_hd__o221a_1
XPHY_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11688_ _11687_/X _11401_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12386_/D sky130_fd_sc_hd__mux2_1
XFILLER_197_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10639_ _11903_/X _10649_/B vssd1 vssd1 vccd1 vccd1 _10639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12309_ _12976_/CLK _12309_/D vssd1 vssd1 vccd1 vccd1 _12309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07850_ _13010_/Q vssd1 vssd1 vccd1 vccd1 _07850_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06801_ _06797_/X _06798_/X _06791_/X _06783_/X _06800_/X vssd1 vssd1 vccd1 vccd1
+ _06801_/X sky130_fd_sc_hd__o221a_1
XFILLER_96_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07781_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07781_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_1
XFILLER_7_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09520_ _09500_/Y _09502_/X _09514_/A vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__o21ai_2
X_06732_ _12026_/X _12023_/X _12029_/X _06731_/X vssd1 vssd1 vccd1 vccd1 _06734_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09451_ _09451_/A vssd1 vssd1 vccd1 vccd1 _09451_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06663_ _06886_/A vssd1 vssd1 vccd1 vccd1 _06663_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_188_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08402_ _08402_/A vssd1 vssd1 vccd1 vccd1 _08418_/A sky130_fd_sc_hd__inv_2
XFILLER_91_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09382_ _09372_/X _09382_/B _09382_/C _09382_/D vssd1 vssd1 vccd1 vccd1 _09382_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_52_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06594_ _06594_/A vssd1 vssd1 vccd1 vccd1 _06598_/A sky130_fd_sc_hd__inv_2
XFILLER_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08333_ _12813_/Q _11588_/X _08335_/S vssd1 vssd1 vccd1 vccd1 _12813_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08264_ _08282_/A vssd1 vssd1 vccd1 vccd1 _08264_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07215_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07215_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_193_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08195_ _13086_/Q _10415_/A _13086_/Q _10415_/A vssd1 vssd1 vccd1 vccd1 _08195_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_192_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07146_ _07161_/A vssd1 vssd1 vccd1 vccd1 _07146_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07077_ _07069_/X _07074_/X _06342_/Y _13149_/Q _07042_/A vssd1 vssd1 vccd1 vccd1
+ _13149_/D sky130_fd_sc_hd__a32o_1
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06028_ _12745_/Q _12713_/Q _06026_/Y _06027_/Y vssd1 vssd1 vccd1 vccd1 _06030_/A
+ sky130_fd_sc_hd__a22o_1
Xoutput373 _11159_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_120_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput384 _11169_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput395 _11179_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__clkbuf_2
XFILLER_75_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07979_ _07985_/A vssd1 vssd1 vccd1 vccd1 _07979_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_132_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09718_ _09747_/A _09825_/A vssd1 vssd1 vccd1 vccd1 _09718_/X sky130_fd_sc_hd__or2_1
XFILLER_142_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10990_ _12539_/Q _12351_/Q _10989_/X vssd1 vssd1 vccd1 vccd1 _10990_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09649_ _12875_/Q vssd1 vssd1 vccd1 vccd1 _09649_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12664_/CLK _12660_/D _08821_/X vssd1 vssd1 vccd1 vccd1 _12660_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11611_ _12493_/Q _12978_/Q _12601_/Q vssd1 vssd1 vccd1 vccd1 _11611_/X sky130_fd_sc_hd__mux2_1
XPHY_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12937_/CLK _12591_/D vssd1 vssd1 vccd1 vccd1 _12591_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ _12831_/Q _10794_/C _11543_/S vssd1 vssd1 vccd1 vccd1 _11542_/X sky130_fd_sc_hd__mux2_1
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11473_ _12916_/Q _09179_/C _11481_/S vssd1 vssd1 vccd1 vccd1 _11473_/X sky130_fd_sc_hd__mux2_1
XPHY_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13212_ _13213_/CLK _13212_/D _06662_/X vssd1 vssd1 vccd1 vccd1 _13212_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10424_ _10429_/C vssd1 vssd1 vccd1 vccd1 _10424_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13143_ _12168_/X _13143_/D _07120_/X vssd1 vssd1 vccd1 vccd1 _13143_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10355_ _10371_/A _10355_/B _10355_/C vssd1 vssd1 vccd1 vccd1 _10355_/Y sky130_fd_sc_hd__nor3_1
XFILLER_140_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10286_ _13160_/Q vssd1 vssd1 vccd1 vccd1 _10286_/Y sky130_fd_sc_hd__inv_2
X_13074_ _12169_/A0 _13074_/D _07311_/X vssd1 vssd1 vccd1 vccd1 _13074_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_151_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12025_ _11085_/X _11076_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _12025_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12927_ _12993_/CLK _12927_/D vssd1 vssd1 vccd1 vccd1 _12927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12858_ _13257_/CLK _12858_/D _08073_/X vssd1 vssd1 vccd1 vccd1 _12858_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_61_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ _09180_/A _11808_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11809_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12166_/A0 _12789_/D _08393_/X vssd1 vssd1 vccd1 vccd1 _12789_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07000_ _11407_/X vssd1 vssd1 vccd1 vccd1 _07012_/A sky130_fd_sc_hd__inv_2
XFILLER_128_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08951_ _12440_/Q _12439_/Q vssd1 vssd1 vccd1 vccd1 _08952_/B sky130_fd_sc_hd__or2_1
XFILLER_102_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07902_ _12920_/Q _11509_/X _07904_/S vssd1 vssd1 vccd1 vccd1 _12920_/D sky130_fd_sc_hd__mux2_1
X_08882_ _08882_/A vssd1 vssd1 vccd1 vccd1 _08882_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07833_ _13031_/Q vssd1 vssd1 vccd1 vccd1 _07833_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07764_ _12590_/Q _07764_/B vssd1 vssd1 vccd1 vccd1 _07765_/B sky130_fd_sc_hd__or2_1
XFILLER_38_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09503_ _09502_/A _09502_/B _09502_/X vssd1 vssd1 vccd1 vccd1 _09504_/B sky130_fd_sc_hd__o21ba_1
X_06715_ _06720_/A _06720_/B vssd1 vssd1 vccd1 vccd1 _06715_/X sky130_fd_sc_hd__or2_1
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07695_ _09268_/B vssd1 vssd1 vccd1 vccd1 _07695_/X sky130_fd_sc_hd__buf_2
X_09434_ _09434_/A _09434_/B _09434_/C vssd1 vssd1 vccd1 vccd1 _09434_/X sky130_fd_sc_hd__or3_2
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06646_ _06886_/A vssd1 vssd1 vccd1 vccd1 _06646_/X sky130_fd_sc_hd__clkbuf_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09365_ _12460_/Q _09356_/Y _09362_/Y _12398_/Q _09364_/X vssd1 vssd1 vccd1 vccd1
+ _09371_/C sky130_fd_sc_hd__o221a_1
XFILLER_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06577_ _13221_/Q vssd1 vssd1 vccd1 vccd1 _06577_/Y sky130_fd_sc_hd__inv_2
X_08316_ _08325_/A vssd1 vssd1 vccd1 vccd1 _08316_/X sky130_fd_sc_hd__clkbuf_1
X_09296_ _09296_/A _09296_/B vssd1 vssd1 vccd1 vccd1 _09296_/X sky130_fd_sc_hd__or2_1
XFILLER_177_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08247_ _08247_/A _08247_/B _08247_/C _08246_/X vssd1 vssd1 vccd1 vccd1 _08275_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_165_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08178_ _13116_/Q _08177_/Y _13139_/Q _08154_/Y vssd1 vssd1 vccd1 vccd1 _08178_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07129_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07129_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10140_ _10140_/A vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10071_ _08272_/Y _10796_/A _08141_/Y _10047_/B vssd1 vssd1 vccd1 vccd1 _10071_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_88_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10973_ _10976_/B _10972_/X _10976_/B _10972_/X vssd1 vssd1 vccd1 vccd1 _12349_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12712_ _12713_/CLK _12712_/D _08674_/X vssd1 vssd1 vccd1 vccd1 _12712_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12643_ _12870_/CLK _12643_/D _08862_/X vssd1 vssd1 vccd1 vccd1 _12643_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12574_ _12976_/CLK _12574_/D vssd1 vssd1 vccd1 vccd1 _12574_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11525_ _12814_/Q _09243_/C _11533_/S vssd1 vssd1 vccd1 vccd1 _11525_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11456_ _12899_/Q input357/X _11459_/S vssd1 vssd1 vccd1 vccd1 _11456_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10407_ _10459_/A vssd1 vssd1 vccd1 vccd1 _10407_/X sky130_fd_sc_hd__buf_2
XFILLER_178_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11387_ _10581_/Y _12401_/D _11392_/S vssd1 vssd1 vccd1 vccd1 _11387_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13126_ _12168_/X _13126_/D _07163_/X vssd1 vssd1 vccd1 vccd1 _13126_/Q sky130_fd_sc_hd__dfrtp_1
X_10338_ _12901_/Q vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__inv_2
XFILLER_140_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_119_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 _12683_/CLK sky130_fd_sc_hd__clkbuf_16
X_13057_ _12165_/X _13057_/D _07363_/X vssd1 vssd1 vccd1 vccd1 _13057_/Q sky130_fd_sc_hd__dfrtp_4
X_10269_ _12634_/Q vssd1 vssd1 vccd1 vccd1 _10269_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12008_ _11114_/X _10737_/X _12193_/S vssd1 vssd1 vccd1 vccd1 _12008_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06500_ _06500_/A _06500_/B vssd1 vssd1 vccd1 vccd1 _06500_/Y sky130_fd_sc_hd__nor2_1
X_07480_ _11456_/X _07474_/X _13015_/Q _07475_/X vssd1 vssd1 vccd1 vccd1 _13015_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06431_ _06356_/X _10738_/A _06427_/X _10737_/A _06430_/X vssd1 vssd1 vccd1 vccd1
+ _06431_/X sky130_fd_sc_hd__o221a_2
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09150_ _09150_/A _12596_/Q _09175_/B vssd1 vssd1 vccd1 vccd1 _09150_/X sky130_fd_sc_hd__or3_4
X_06362_ _13253_/Q vssd1 vssd1 vccd1 vccd1 _06362_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_194_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08101_ _08257_/A vssd1 vssd1 vccd1 vccd1 _08101_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09081_ _12546_/Q _09079_/A _09180_/B _09079_/Y vssd1 vssd1 vccd1 vccd1 _12546_/D
+ sky130_fd_sc_hd__a22o_1
X_06293_ _06313_/A vssd1 vssd1 vccd1 vccd1 _06293_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08032_ _08036_/A vssd1 vssd1 vccd1 vccd1 _08032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput50 la_data_in[10] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_1
XFILLER_116_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput61 la_data_in[11] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_1
Xinput72 la_data_in[14] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_1
XFILLER_190_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput83 la_data_in[24] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__buf_1
XFILLER_157_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput94 la_data_in[34] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__buf_1
XFILLER_192_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09983_ _12637_/Q vssd1 vssd1 vccd1 vccd1 _09983_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08934_ _12441_/Q _12442_/Q vssd1 vssd1 vccd1 vccd1 _11916_/S sky130_fd_sc_hd__nor2_1
XFILLER_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08865_ _07747_/X _06332_/Y _08852_/X _12642_/Q vssd1 vssd1 vccd1 vccd1 _12642_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater640 input341/X vssd1 vssd1 vccd1 vccd1 _09180_/B sky130_fd_sc_hd__buf_8
Xrepeater651 _07993_/A vssd1 vssd1 vccd1 vccd1 _09243_/C sky130_fd_sc_hd__buf_8
X_07816_ _13018_/Q vssd1 vssd1 vccd1 vccd1 _07816_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08796_ _08807_/A vssd1 vssd1 vccd1 vccd1 _08796_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07747_ _08849_/A vssd1 vssd1 vccd1 vccd1 _07747_/X sky130_fd_sc_hd__buf_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07678_ _07678_/A _07678_/B _07678_/C vssd1 vssd1 vccd1 vccd1 _07685_/A sky130_fd_sc_hd__nor3_4
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09417_ _12452_/Q _09390_/Y _12458_/Q _09385_/Y _09416_/X vssd1 vssd1 vccd1 vccd1
+ _09422_/C sky130_fd_sc_hd__a221o_1
X_06629_ _06650_/A vssd1 vssd1 vccd1 vccd1 _06629_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_179_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09348_ _12542_/Q _09346_/Y _09338_/Y _12409_/Q _09347_/X vssd1 vssd1 vccd1 vccd1
+ _09353_/C sky130_fd_sc_hd__o221a_1
XFILLER_12_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _09279_/A _09279_/B _09279_/C _09279_/D vssd1 vssd1 vccd1 vccd1 _09279_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ vssd1 vssd1 vccd1 vccd1 _11310_/HI _11310_/LO sky130_fd_sc_hd__conb_1
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12290_ _12296_/CLK _12290_/D vssd1 vssd1 vccd1 vccd1 _12290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11241_ vssd1 vssd1 vccd1 vccd1 _11241_/HI _11241_/LO sky130_fd_sc_hd__conb_1
XFILLER_107_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11172_ vssd1 vssd1 vccd1 vccd1 _11172_/HI _11172_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10123_ _13259_/Q vssd1 vssd1 vccd1 vccd1 _10123_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10054_ _10054_/A _10796_/A vssd1 vssd1 vccd1 vccd1 _10054_/Y sky130_fd_sc_hd__nor2_2
XFILLER_76_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10956_ _12535_/Q vssd1 vssd1 vccd1 vccd1 _10958_/A sky130_fd_sc_hd__inv_2
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10887_ _10888_/D _10886_/X _10888_/D _10886_/X vssd1 vssd1 vccd1 vccd1 _12337_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ _12646_/CLK _12626_/D _08905_/X vssd1 vssd1 vccd1 vccd1 _12626_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12557_ _12558_/CLK _12557_/D vssd1 vssd1 vccd1 vccd1 _12557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11508_ _10389_/X _10794_/D _11513_/S vssd1 vssd1 vccd1 vccd1 _11508_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12488_ _12489_/CLK _12488_/D vssd1 vssd1 vccd1 vccd1 _12488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11439_ _12914_/Q _09180_/A _11443_/S vssd1 vssd1 vccd1 vccd1 _11439_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13109_ _12167_/X _13109_/D _07213_/X vssd1 vssd1 vccd1 vccd1 _13109_/Q sky130_fd_sc_hd__dfrtp_1
X_06980_ _06980_/A vssd1 vssd1 vccd1 vccd1 _13177_/D sky130_fd_sc_hd__inv_2
XFILLER_113_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08650_ _11930_/X _08639_/X _12721_/Q _08640_/X vssd1 vssd1 vccd1 vccd1 _12721_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07601_ _12976_/Q _07600_/B _07599_/Y _07600_/Y vssd1 vssd1 vccd1 vccd1 _07602_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08581_ _08591_/A vssd1 vssd1 vccd1 vccd1 _08581_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_87_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _12765_/CLK sky130_fd_sc_hd__clkbuf_16
X_07532_ _07532_/A vssd1 vssd1 vccd1 vccd1 _07532_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_16_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12168_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07463_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07463_/X sky130_fd_sc_hd__clkbuf_1
X_09202_ _12485_/Q _09199_/X _09179_/B _09200_/X vssd1 vssd1 vccd1 vccd1 _12485_/D
+ sky130_fd_sc_hd__a22o_1
X_06414_ _06887_/A vssd1 vssd1 vccd1 vccd1 _06415_/B sky130_fd_sc_hd__clkbuf_2
X_07394_ _07408_/A vssd1 vssd1 vccd1 vccd1 _07394_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09133_ _12306_/Q vssd1 vssd1 vccd1 vccd1 _09152_/A sky130_fd_sc_hd__inv_2
XFILLER_33_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06345_ _06122_/A _06122_/B _06122_/Y vssd1 vssd1 vccd1 vccd1 _06346_/A sky130_fd_sc_hd__o21ai_4
XFILLER_175_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06276_ _06072_/Y _06073_/Y _06075_/B _06181_/X vssd1 vssd1 vccd1 vccd1 _06276_/X
+ sky130_fd_sc_hd__o22a_1
X_09064_ _09067_/A vssd1 vssd1 vccd1 vccd1 _09064_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08015_ _12879_/Q _07996_/A _07304_/X _07998_/A vssd1 vssd1 vccd1 vccd1 _12879_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09966_ _10034_/A _10113_/A vssd1 vssd1 vccd1 vccd1 _10010_/A sky130_fd_sc_hd__or2_2
XFILLER_44_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08917_ _08962_/A vssd1 vssd1 vccd1 vccd1 _08917_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09897_ _09897_/A vssd1 vssd1 vccd1 vccd1 _09897_/X sky130_fd_sc_hd__buf_2
XFILLER_100_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08848_ _08851_/A vssd1 vssd1 vccd1 vccd1 _08848_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08779_ _08789_/A vssd1 vssd1 vccd1 vccd1 _08779_/X sky130_fd_sc_hd__clkbuf_1
XPHY_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _12513_/Q _12325_/Q vssd1 vssd1 vccd1 vccd1 _10810_/Y sky130_fd_sc_hd__nor2_1
XPHY_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11789_/X _12130_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12437_/D sky130_fd_sc_hd__mux2_1
XPHY_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10741_ _13251_/Q vssd1 vssd1 vccd1 vccd1 _10742_/A sky130_fd_sc_hd__inv_2
XPHY_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10672_ _12433_/Q _12434_/Q _12435_/Q vssd1 vssd1 vccd1 vccd1 _10672_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12411_ _12547_/CLK _12411_/D vssd1 vssd1 vccd1 vccd1 _12411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12342_ _12529_/CLK _12342_/D vssd1 vssd1 vccd1 vccd1 _12342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12273_ _10176_/X _12899_/Q _11867_/X _11868_/X _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12289_/D sky130_fd_sc_hd__mux4_2
XFILLER_5_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11224_ vssd1 vssd1 vccd1 vccd1 _11224_/HI _11224_/LO sky130_fd_sc_hd__conb_1
XFILLER_153_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11155_ vssd1 vssd1 vccd1 vccd1 _11155_/HI _11155_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10106_ _10103_/Y _09999_/A _09507_/Y _10141_/A _10105_/X vssd1 vssd1 vccd1 vccd1
+ _10107_/D sky130_fd_sc_hd__o221a_1
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11086_ _11086_/A vssd1 vssd1 vccd1 vccd1 _11086_/X sky130_fd_sc_hd__clkbuf_2
Xinput240 la_oenb[50] vssd1 vssd1 vccd1 vccd1 input240/X sky130_fd_sc_hd__buf_1
XFILLER_88_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput251 la_oenb[60] vssd1 vssd1 vccd1 vccd1 input251/X sky130_fd_sc_hd__buf_1
XFILLER_0_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput262 la_oenb[70] vssd1 vssd1 vccd1 vccd1 input262/X sky130_fd_sc_hd__buf_1
X_10037_ _12772_/Q vssd1 vssd1 vccd1 vccd1 _10037_/Y sky130_fd_sc_hd__inv_2
Xinput273 la_oenb[80] vssd1 vssd1 vccd1 vccd1 input273/X sky130_fd_sc_hd__buf_1
Xinput284 la_oenb[90] vssd1 vssd1 vccd1 vccd1 input284/X sky130_fd_sc_hd__buf_1
XFILLER_64_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput295 wb_rst_i vssd1 vssd1 vccd1 vccd1 _07590_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_64_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11988_ _11127_/X _11120_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10939_ _12531_/Q _12343_/Q _10930_/Y _10933_/Y vssd1 vssd1 vccd1 vccd1 _10939_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _13268_/CLK _12610_/Q _08969_/X vssd1 vssd1 vccd1 vccd1 _12609_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06130_ _06130_/A _06130_/B _06130_/C vssd1 vssd1 vccd1 vccd1 _06130_/X sky130_fd_sc_hd__and3_1
XFILLER_200_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_134_wb_clk_i _12726_/CLK vssd1 vssd1 vccd1 vccd1 _13161_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06061_ _12733_/Q _12701_/Q vssd1 vssd1 vccd1 vccd1 _06064_/A sky130_fd_sc_hd__nand2_2
XFILLER_144_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09820_ _06529_/Y _06533_/Y _09810_/Y _09812_/Y vssd1 vssd1 vccd1 vccd1 _09820_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09751_ _09751_/A _09751_/B vssd1 vssd1 vccd1 vccd1 _09849_/A sky130_fd_sc_hd__nand2_2
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06963_ _11854_/X _06960_/B _06961_/B vssd1 vssd1 vccd1 vccd1 _06963_/X sky130_fd_sc_hd__a21bo_1
X_08702_ _11835_/X _08700_/X _12701_/Q _08701_/X vssd1 vssd1 vccd1 vccd1 _12701_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09682_ _09886_/A vssd1 vssd1 vccd1 vccd1 _09682_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06894_ _06916_/A vssd1 vssd1 vccd1 vccd1 _06894_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08633_ _11937_/X _08624_/X _12728_/Q _08625_/X vssd1 vssd1 vccd1 vccd1 _12728_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _08817_/A vssd1 vssd1 vccd1 vccd1 _08781_/A sky130_fd_sc_hd__buf_2
XFILLER_70_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07515_ _07515_/A vssd1 vssd1 vccd1 vccd1 _10527_/B sky130_fd_sc_hd__clkbuf_4
XPHY_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08495_ _12771_/Q _08494_/X _09019_/A _07888_/A vssd1 vssd1 vccd1 vccd1 _12771_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07446_ _11469_/X _07444_/X _13028_/Q _07445_/X vssd1 vssd1 vccd1 vccd1 _13028_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07377_ _07477_/A vssd1 vssd1 vccd1 vccd1 _07462_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09116_ _09116_/A vssd1 vssd1 vccd1 vccd1 _09116_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06328_ _06303_/X _06314_/X _06327_/Y _13260_/Q _06306_/X vssd1 vssd1 vccd1 vccd1
+ _13260_/D sky130_fd_sc_hd__a32o_1
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09047_ _09051_/A _12158_/X vssd1 vssd1 vccd1 vccd1 _12569_/D sky130_fd_sc_hd__nor2b_1
XFILLER_50_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06259_ _06259_/A vssd1 vssd1 vccd1 vccd1 _06259_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09949_ _09949_/A vssd1 vssd1 vccd1 vccd1 _09949_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12960_ _12960_/CLK _12960_/D vssd1 vssd1 vccd1 vccd1 _12960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11911_ _12441_/Q _11910_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _11911_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12891_ _12892_/CLK _12891_/D _07979_/X vssd1 vssd1 vccd1 vccd1 _12891_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _09953_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11842_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _12115_/X _11772_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11773_/X sky130_fd_sc_hd__mux2_1
XPHY_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _13249_/Q vssd1 vssd1 vccd1 vccd1 _10758_/A sky130_fd_sc_hd__inv_2
XFILLER_198_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10655_ _11909_/X _10655_/B vssd1 vssd1 vccd1 vccd1 _10655_/X sky130_fd_sc_hd__and2_1
XFILLER_186_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10586_ _10586_/A _10586_/B vssd1 vssd1 vccd1 vccd1 _10594_/A sky130_fd_sc_hd__nor2_4
XFILLER_6_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12325_ _12999_/CLK _12325_/D vssd1 vssd1 vccd1 vccd1 _12325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12256_ _12255_/X _12648_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12256_/X sky130_fd_sc_hd__mux2_2
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_11207_ vssd1 vssd1 vccd1 vccd1 _11207_/HI _11207_/LO sky130_fd_sc_hd__conb_1
XFILLER_141_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12187_ _11062_/A _11049_/A _12200_/S vssd1 vssd1 vccd1 vccd1 _12187_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11138_ _10763_/A _10788_/A _13248_/Q _11111_/X _11112_/X vssd1 vssd1 vccd1 vccd1
+ _11138_/X sky130_fd_sc_hd__a221o_1
XFILLER_122_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11069_ _10693_/X _10759_/X _06407_/X _10760_/X _10761_/X vssd1 vssd1 vccd1 vccd1
+ _11069_/X sky130_fd_sc_hd__a221o_1
XFILLER_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07300_ _07562_/A vssd1 vssd1 vccd1 vccd1 _07300_/X sky130_fd_sc_hd__buf_2
X_08280_ _08353_/S vssd1 vssd1 vccd1 vccd1 _08292_/S sky130_fd_sc_hd__buf_2
XFILLER_20_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07231_ _11567_/X _07218_/X _13102_/Q _07219_/X vssd1 vssd1 vccd1 vccd1 _13102_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07162_ _11528_/X _07160_/X _13127_/Q _07161_/X vssd1 vssd1 vccd1 vccd1 _13127_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06113_ _12689_/Q vssd1 vssd1 vccd1 vccd1 _06113_/Y sky130_fd_sc_hd__inv_2
X_07093_ _09267_/B vssd1 vssd1 vccd1 vccd1 _09071_/A sky130_fd_sc_hd__inv_2
XFILLER_145_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput500 _11249_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_201_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput511 _11259_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput522 _11269_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__clkbuf_2
X_06044_ _12742_/Q _12710_/Q _12742_/Q _12710_/Q vssd1 vssd1 vccd1 vccd1 _06044_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
Xoutput533 _11279_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__clkbuf_2
Xoutput544 _11289_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput555 _11299_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__clkbuf_2
Xoutput566 _11309_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput577 _12294_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput588 _12560_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput599 _12570_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09803_ _09803_/A _09824_/A vssd1 vssd1 vccd1 vccd1 _09803_/X sky130_fd_sc_hd__or2_1
XFILLER_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07995_ _08004_/A vssd1 vssd1 vccd1 vccd1 _07995_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09734_ _09731_/Y _09733_/A _09747_/B _09733_/Y _09701_/A vssd1 vssd1 vccd1 vccd1
+ _09735_/B sky130_fd_sc_hd__o221a_1
XFILLER_189_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06946_ _12055_/X _06944_/Y _12054_/X _06945_/X vssd1 vssd1 vccd1 vccd1 _06946_/X
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12426_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ _13200_/Q vssd1 vssd1 vccd1 vccd1 _09665_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06877_ _06874_/X _06875_/X _12000_/X _06876_/X vssd1 vssd1 vccd1 vccd1 _06877_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08616_ _11944_/X _08608_/X _12735_/Q _08610_/X vssd1 vssd1 vccd1 vccd1 _12735_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09596_ _09595_/Y _07735_/A _12871_/Q _12614_/Q vssd1 vssd1 vccd1 vccd1 _09596_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _07737_/A _07059_/A _12045_/X _08546_/Y _07074_/X vssd1 vssd1 vccd1 vccd1
+ _08548_/A sky130_fd_sc_hd__o32a_1
XPHY_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08478_ _13071_/Q _10395_/A _13055_/Q _10352_/A vssd1 vssd1 vccd1 vccd1 _08478_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07429_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07429_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10440_ _10444_/C vssd1 vssd1 vccd1 vccd1 _10442_/B sky130_fd_sc_hd__inv_2
XFILLER_148_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10371_ _10371_/A _10376_/C _10371_/C vssd1 vssd1 vccd1 vccd1 _10371_/Y sky130_fd_sc_hd__nor3_1
XFILLER_3_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12110_ _12109_/X _12432_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12110_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13090_ _12167_/X _13090_/D _07260_/X vssd1 vssd1 vccd1 vccd1 _13090_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12041_ _10791_/X _10790_/Y _12193_/S vssd1 vssd1 vccd1 vccd1 _12041_/X sky130_fd_sc_hd__mux2_2
XFILLER_123_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12943_ _13260_/CLK _12943_/D _07739_/X vssd1 vssd1 vccd1 vccd1 _12943_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12874_ _12875_/CLK _12874_/D _08030_/X vssd1 vssd1 vccd1 vccd1 _12874_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _09908_/Y _12850_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11825_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11756_ _09186_/A _11755_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11756_/X sky130_fd_sc_hd__mux2_1
XPHY_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _12765_/Q _12764_/Q vssd1 vssd1 vccd1 vccd1 _10707_/Y sky130_fd_sc_hd__nor2_2
XPHY_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11687_ _11401_/X _10528_/C _11691_/S vssd1 vssd1 vccd1 vccd1 _11687_/X sky130_fd_sc_hd__mux2_1
XPHY_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10638_ _11903_/X vssd1 vssd1 vccd1 vccd1 _10638_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10569_ _10521_/A _09411_/Y _09423_/Y _12395_/D _10562_/A vssd1 vssd1 vccd1 vccd1
+ _10570_/B sky130_fd_sc_hd__o32a_1
XFILLER_6_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12308_ _12976_/CLK _12308_/D vssd1 vssd1 vccd1 vccd1 _12308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12239_ _12774_/Q _12847_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12239_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06800_ _10717_/A _06804_/B vssd1 vssd1 vccd1 vccd1 _06800_/X sky130_fd_sc_hd__or2_1
XFILLER_7_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07780_ _07780_/A vssd1 vssd1 vccd1 vccd1 _07780_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_1
XFILLER_77_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06731_ _12026_/X _12023_/X _12026_/X _12023_/X vssd1 vssd1 vccd1 vccd1 _06731_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09450_ _12928_/Q _09438_/X _13004_/Q _09442_/X vssd1 vssd1 vccd1 vccd1 _09450_/X
+ sky130_fd_sc_hd__a22o_1
X_06662_ _06690_/A vssd1 vssd1 vccd1 vccd1 _06662_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08401_ _08417_/A vssd1 vssd1 vccd1 vccd1 _08401_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_197_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09381_ _12454_/Q _09367_/Y _12459_/Q _09337_/Y _09380_/X vssd1 vssd1 vccd1 vccd1
+ _09382_/D sky130_fd_sc_hd__o221a_1
XFILLER_36_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06593_ _12202_/X _12201_/X _06587_/X _06588_/X _06592_/X vssd1 vssd1 vccd1 vccd1
+ _06594_/A sky130_fd_sc_hd__o32a_1
XFILLER_149_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08332_ _08339_/A vssd1 vssd1 vccd1 vccd1 _08332_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08263_ _12838_/Q _08251_/X _07304_/X _11417_/S vssd1 vssd1 vccd1 vccd1 _12838_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07214_ _11574_/X _07201_/X _13109_/Q _07204_/X vssd1 vssd1 vccd1 vccd1 _13109_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08194_ _13084_/Q vssd1 vssd1 vccd1 vccd1 _08194_/Y sky130_fd_sc_hd__inv_2
X_07145_ _07160_/A vssd1 vssd1 vccd1 vccd1 _07145_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07076_ _07078_/A vssd1 vssd1 vccd1 vccd1 _07076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06027_ _12713_/Q vssd1 vssd1 vccd1 vccd1 _06027_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput374 _11160_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput385 _11170_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__clkbuf_2
Xoutput396 _11180_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07978_ _12892_/Q _07974_/X _07975_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _12892_/D
+ sky130_fd_sc_hd__a22o_1
X_09717_ _09717_/A _09717_/B vssd1 vssd1 vccd1 vccd1 _09825_/A sky130_fd_sc_hd__nand2_2
XFILLER_68_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06929_ _06926_/X _06927_/X _12005_/X _06928_/X vssd1 vssd1 vccd1 vccd1 _06929_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09648_ _13160_/Q _09475_/X _09629_/Y _09919_/B _09647_/X vssd1 vssd1 vccd1 vccd1
+ _09648_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09578_/A _09578_/B _09578_/C vssd1 vssd1 vccd1 vccd1 _09580_/B sky130_fd_sc_hd__o21a_1
XFILLER_169_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _10487_/X _10793_/A _11610_/S vssd1 vssd1 vccd1 vccd1 _11610_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12937_/CLK _12590_/D vssd1 vssd1 vccd1 vccd1 _12590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _12830_/Q _10794_/D _11543_/S vssd1 vssd1 vccd1 vccd1 _11541_/X sky130_fd_sc_hd__mux2_1
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ _12915_/Q _09179_/D _11481_/S vssd1 vssd1 vccd1 vccd1 _11472_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13211_ _13213_/CLK _13211_/D _06676_/X vssd1 vssd1 vccd1 vccd1 _13211_/Q sky130_fd_sc_hd__dfrtp_1
X_10423_ _08117_/X _10422_/B _10429_/C _10407_/X vssd1 vssd1 vccd1 vccd1 _10423_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13142_ _12168_/X _13142_/D _07122_/X vssd1 vssd1 vccd1 vccd1 _13142_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10354_ _07839_/X _10352_/C _10352_/A vssd1 vssd1 vccd1 vccd1 _10355_/C sky130_fd_sc_hd__o21a_1
XFILLER_87_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13073_ _12165_/X _13073_/D _07315_/X vssd1 vssd1 vccd1 vccd1 _13073_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10285_ _12635_/Q vssd1 vssd1 vccd1 vccd1 _10285_/Y sky130_fd_sc_hd__inv_2
X_12024_ _11068_/X _11063_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _12024_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12926_ _12993_/CLK _12926_/D vssd1 vssd1 vccd1 vccd1 _12926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12857_ _13257_/CLK _12857_/D _08075_/X vssd1 vssd1 vccd1 vccd1 _12857_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _12079_/X _12490_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__mux2_1
X_12788_ _12872_/CLK _12788_/D _08395_/X vssd1 vssd1 vccd1 vccd1 _12788_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11739_ _11369_/X _12469_/Q _12103_/S vssd1 vssd1 vccd1 vccd1 _11739_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08950_ _12437_/Q _12438_/Q vssd1 vssd1 vccd1 vccd1 _09315_/A sky130_fd_sc_hd__or2_2
XFILLER_143_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07901_ _07903_/A vssd1 vssd1 vccd1 vccd1 _07901_/X sky130_fd_sc_hd__clkbuf_1
X_08881_ _08877_/X _06278_/Y _08878_/X _12636_/Q vssd1 vssd1 vccd1 vccd1 _12636_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_29_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07832_ _12923_/Q vssd1 vssd1 vccd1 vccd1 _10397_/A sky130_fd_sc_hd__buf_2
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07763_ _12589_/Q _07763_/B vssd1 vssd1 vccd1 vccd1 _07764_/B sky130_fd_sc_hd__or2_1
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09502_ _09502_/A _09502_/B vssd1 vssd1 vccd1 vccd1 _09502_/X sky130_fd_sc_hd__and2_1
X_06714_ _06711_/X _06712_/X _06711_/X _06712_/X vssd1 vssd1 vccd1 vccd1 _06720_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07694_ _07717_/A vssd1 vssd1 vccd1 vccd1 _07694_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09433_ _09433_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09434_/C sky130_fd_sc_hd__nor2_1
X_06645_ _11901_/X _12196_/X _06639_/X _06640_/X _06644_/X vssd1 vssd1 vccd1 vccd1
+ _06645_/X sky130_fd_sc_hd__o32a_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _09335_/Y _12397_/Q _09363_/Y _12414_/Q vssd1 vssd1 vccd1 vccd1 _09364_/X
+ sky130_fd_sc_hd__o22a_1
X_06576_ _06576_/A _06576_/B vssd1 vssd1 vccd1 vccd1 _06576_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08315_ _12821_/Q _11596_/X _08321_/S vssd1 vssd1 vccd1 vccd1 _12821_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09295_ _09295_/A _09296_/B vssd1 vssd1 vccd1 vccd1 _11348_/S sky130_fd_sc_hd__or2_4
XFILLER_177_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08246_ _08240_/X _08246_/B _08246_/C _08246_/D vssd1 vssd1 vccd1 vccd1 _08246_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_123_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08177_ _12806_/Q vssd1 vssd1 vccd1 vccd1 _08177_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07128_ _11541_/X _07113_/X _13140_/Q _07116_/X vssd1 vssd1 vccd1 vccd1 _13140_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07059_ _07059_/A vssd1 vssd1 vccd1 vccd1 _07059_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10070_ _10151_/A vssd1 vssd1 vccd1 vccd1 _10070_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10972_ _10962_/Y _10963_/Y _10976_/A _10967_/X vssd1 vssd1 vccd1 vccd1 _10972_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_29_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ _12713_/CLK _12711_/D _08676_/X vssd1 vssd1 vccd1 vccd1 _12711_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_71_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ _12870_/CLK _12642_/D _08864_/X vssd1 vssd1 vccd1 vccd1 _12642_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12573_ _12976_/CLK _12573_/D vssd1 vssd1 vccd1 vccd1 _12573_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11524_ _12813_/Q _09243_/D _11533_/S vssd1 vssd1 vccd1 vccd1 _11524_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11455_ _12898_/Q input356/X _11459_/S vssd1 vssd1 vccd1 vccd1 _11455_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10406_ _10411_/A vssd1 vssd1 vccd1 vccd1 _10459_/A sky130_fd_sc_hd__inv_2
XFILLER_109_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11386_ _10582_/X _12402_/D _11390_/S vssd1 vssd1 vccd1 vccd1 _11386_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13125_ _12168_/X _13125_/D _07165_/X vssd1 vssd1 vccd1 vccd1 _13125_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10337_ _10342_/C vssd1 vssd1 vccd1 vccd1 _10337_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13056_ _12165_/X _13056_/D _07365_/X vssd1 vssd1 vccd1 vccd1 _13056_/Q sky130_fd_sc_hd__dfrtp_4
X_10268_ _12889_/Q vssd1 vssd1 vccd1 vccd1 _10268_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12007_ _11113_/X _11110_/Y _12199_/S vssd1 vssd1 vccd1 vccd1 _12007_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10199_ _12869_/Q vssd1 vssd1 vccd1 vccd1 _10199_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_159_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12537_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12909_ _12166_/X _12909_/D _07927_/X vssd1 vssd1 vccd1 vccd1 _12909_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06430_ _06430_/A vssd1 vssd1 vccd1 vccd1 _06430_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06361_ _08504_/A vssd1 vssd1 vccd1 vccd1 _06361_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_187_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08100_ _08284_/A vssd1 vssd1 vccd1 vccd1 _08257_/A sky130_fd_sc_hd__clkbuf_2
X_09080_ _12547_/Q _09079_/A _09180_/A _09079_/Y vssd1 vssd1 vccd1 vccd1 _12547_/D
+ sky130_fd_sc_hd__a22o_1
X_06292_ _06269_/X _06281_/X _06291_/Y _13267_/Q _06273_/X vssd1 vssd1 vccd1 vccd1
+ _13267_/D sky130_fd_sc_hd__a32o_1
X_08031_ _12874_/Q _08024_/X _07983_/X _08026_/X vssd1 vssd1 vccd1 vccd1 _12874_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput40 la_data_in[100] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_1
Xinput51 la_data_in[110] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_1
Xinput62 la_data_in[120] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_1
Xinput73 la_data_in[15] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_1
Xinput84 la_data_in[25] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__buf_1
XFILLER_196_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput95 la_data_in[35] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__buf_1
XFILLER_190_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09982_ _09984_/A _09982_/B _11967_/S _09982_/D vssd1 vssd1 vccd1 vccd1 _10166_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08933_ _12444_/Q vssd1 vssd1 vccd1 vccd1 _08936_/A sky130_fd_sc_hd__inv_2
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08864_ _08866_/A vssd1 vssd1 vccd1 vccd1 _08864_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater630 _11522_/S vssd1 vssd1 vccd1 vccd1 _11546_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_84_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07815_ _12914_/Q vssd1 vssd1 vccd1 vccd1 _07815_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater641 input340/X vssd1 vssd1 vccd1 vccd1 _09185_/D sky130_fd_sc_hd__buf_8
Xrepeater652 input329/X vssd1 vssd1 vccd1 vccd1 _09184_/A sky130_fd_sc_hd__buf_8
X_08795_ _08794_/Y _08781_/X _06265_/X _08764_/A vssd1 vssd1 vccd1 vccd1 _12670_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_123_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07746_ _08849_/A vssd1 vssd1 vccd1 vccd1 _07746_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07677_ _12965_/Q _07676_/B _09283_/A _07676_/Y vssd1 vssd1 vccd1 vccd1 _12965_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09416_ _12466_/Q _09415_/Y _12545_/Q _09399_/Y vssd1 vssd1 vccd1 vccd1 _09416_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06628_ _06628_/A vssd1 vssd1 vccd1 vccd1 _13216_/D sky130_fd_sc_hd__inv_2
XFILLER_186_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09347_ _12465_/Q _12401_/Q _12465_/Q _12401_/Q vssd1 vssd1 vccd1 vccd1 _09347_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_166_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06559_ _06559_/A vssd1 vssd1 vccd1 vccd1 _13223_/D sky130_fd_sc_hd__inv_2
XFILLER_179_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09278_ _09278_/A vssd1 vssd1 vccd1 vccd1 _09278_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08229_ _13100_/Q vssd1 vssd1 vccd1 vccd1 _08229_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ vssd1 vssd1 vccd1 vccd1 _11240_/HI _11240_/LO sky130_fd_sc_hd__conb_1
XFILLER_107_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11171_ vssd1 vssd1 vccd1 vccd1 _11171_/HI _11171_/LO sky130_fd_sc_hd__conb_1
XFILLER_84_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10122_ _10121_/Y _10137_/A _09903_/Y _10003_/A vssd1 vssd1 vccd1 vccd1 _10128_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10053_ _13082_/Q _10049_/X _13114_/Q _10051_/X _10052_/Y vssd1 vssd1 vccd1 vccd1
+ _10053_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10955_ _10977_/D _10977_/A _10977_/D _10977_/A vssd1 vssd1 vccd1 vccd1 _12346_/D
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_113_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10886_ _10879_/Y _10880_/Y _10888_/C _10882_/Y vssd1 vssd1 vccd1 vccd1 _10886_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12625_ _12646_/CLK _12625_/D _08907_/X vssd1 vssd1 vccd1 vccd1 _12625_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12556_ _12558_/CLK _12556_/D vssd1 vssd1 vccd1 vccd1 _12556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11507_ _10387_/Y _10792_/A _11513_/S vssd1 vssd1 vccd1 vccd1 _11507_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12487_ _12489_/CLK _12487_/D vssd1 vssd1 vccd1 vccd1 _12487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11438_ _12913_/Q _09180_/B _11443_/S vssd1 vssd1 vccd1 vccd1 _11438_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11369_ _11368_/X _12425_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _11369_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13108_ _12167_/X _13108_/D _07215_/X vssd1 vssd1 vccd1 vccd1 _13108_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13039_ _12164_/X _13039_/D _07418_/X vssd1 vssd1 vccd1 vccd1 _13039_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07600_ _12976_/Q _07600_/B vssd1 vssd1 vccd1 vccd1 _07600_/Y sky130_fd_sc_hd__nand2_1
X_08580_ _08642_/A vssd1 vssd1 vccd1 vccd1 _08591_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07531_ _07531_/A vssd1 vssd1 vccd1 vccd1 _07531_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07462_ _07462_/A vssd1 vssd1 vccd1 vccd1 _07473_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_168_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09201_ _12486_/Q _09199_/X _09179_/A _09200_/X vssd1 vssd1 vccd1 vccd1 _12486_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06413_ _12621_/Q vssd1 vssd1 vccd1 vccd1 _06887_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07393_ _07462_/A vssd1 vssd1 vccd1 vccd1 _07408_/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_56_wb_clk_i _12328_/CLK vssd1 vssd1 vccd1 vccd1 _12773_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09132_ _12510_/Q _09115_/A _07568_/X _09116_/A vssd1 vssd1 vccd1 vccd1 _12510_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06344_ _06344_/A vssd1 vssd1 vccd1 vccd1 _06344_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ _10227_/A _12144_/X vssd1 vssd1 vccd1 vccd1 _12555_/D sky130_fd_sc_hd__nor2b_4
X_06275_ _06280_/A vssd1 vssd1 vccd1 vccd1 _06275_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08014_ _08018_/A vssd1 vssd1 vccd1 vccd1 _08014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09965_ _09981_/A vssd1 vssd1 vccd1 vccd1 _10034_/A sky130_fd_sc_hd__inv_2
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08916_ _08898_/A _06351_/A _08908_/X _12622_/Q vssd1 vssd1 vccd1 vccd1 _12622_/D
+ sky130_fd_sc_hd__o22a_1
X_09896_ _12656_/Q vssd1 vssd1 vccd1 vccd1 _09896_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08847_ _07746_/X _06295_/Y _08837_/X _12649_/Q vssd1 vssd1 vccd1 vccd1 _12649_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08778_ _08777_/Y _08760_/X _06237_/X _08764_/X vssd1 vssd1 vccd1 vccd1 _12675_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _12614_/Q vssd1 vssd1 vccd1 vccd1 _07729_/X sky130_fd_sc_hd__buf_2
XPHY_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _10736_/X _10737_/X _06365_/X _10738_/X _10739_/X vssd1 vssd1 vccd1 vccd1
+ _10740_/X sky130_fd_sc_hd__a221o_1
XPHY_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10671_ _12433_/Q _12434_/Q vssd1 vssd1 vccd1 vccd1 _10671_/X sky130_fd_sc_hd__and2_1
XFILLER_129_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12410_ _12410_/CLK _12410_/D vssd1 vssd1 vccd1 vccd1 _12410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12341_ _12529_/CLK _12341_/D vssd1 vssd1 vccd1 vccd1 _12341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12272_ _10155_/Y _12898_/Q _11865_/X _11866_/X _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12288_/D sky130_fd_sc_hd__mux4_2
XFILLER_182_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11223_ vssd1 vssd1 vccd1 vccd1 _11223_/HI _11223_/LO sky130_fd_sc_hd__conb_1
XFILLER_175_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11154_ vssd1 vssd1 vccd1 vccd1 _11154_/HI _11154_/LO sky130_fd_sc_hd__conb_1
XFILLER_175_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10105_ _10792_/D _10035_/A _08553_/Y _10104_/Y _10140_/A vssd1 vssd1 vccd1 vccd1
+ _10105_/X sky130_fd_sc_hd__o32a_1
XFILLER_89_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11085_ _11041_/X _11075_/X _06392_/X _11083_/X _11084_/X vssd1 vssd1 vccd1 vccd1
+ _11085_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput230 la_oenb[41] vssd1 vssd1 vccd1 vccd1 input230/X sky130_fd_sc_hd__buf_1
Xinput241 la_oenb[51] vssd1 vssd1 vccd1 vccd1 input241/X sky130_fd_sc_hd__buf_1
XFILLER_49_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput252 la_oenb[61] vssd1 vssd1 vccd1 vccd1 input252/X sky130_fd_sc_hd__buf_1
X_10036_ _12754_/Q vssd1 vssd1 vccd1 vccd1 _10036_/Y sky130_fd_sc_hd__inv_2
Xinput263 la_oenb[71] vssd1 vssd1 vccd1 vccd1 input263/X sky130_fd_sc_hd__buf_1
Xinput274 la_oenb[81] vssd1 vssd1 vccd1 vccd1 input274/X sky130_fd_sc_hd__buf_1
Xinput285 la_oenb[91] vssd1 vssd1 vccd1 vccd1 input285/X sky130_fd_sc_hd__buf_1
XFILLER_64_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput296 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _07547_/A sky130_fd_sc_hd__buf_4
XFILLER_5_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ _11124_/X _11117_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _11987_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10938_ _10936_/Y _10937_/Y _12532_/Q _12344_/Q vssd1 vssd1 vccd1 vccd1 _10945_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10869_ _10836_/Y _10864_/X _10890_/C vssd1 vssd1 vccd1 vccd1 _10869_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _13257_/CLK _12609_/Q _08971_/X vssd1 vssd1 vccd1 vccd1 _12608_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12539_ _12540_/CLK _12539_/D vssd1 vssd1 vccd1 vccd1 _12539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06060_ _06060_/A _06259_/A vssd1 vssd1 vccd1 vccd1 _06172_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_103_wb_clk_i _13235_/CLK vssd1 vssd1 vccd1 vccd1 _13227_/CLK sky130_fd_sc_hd__clkbuf_16
X_09750_ _09715_/Y _09770_/A _09749_/Y vssd1 vssd1 vccd1 vccd1 _09751_/B sky130_fd_sc_hd__o21a_1
X_06962_ _11408_/X _11394_/X _06961_/A vssd1 vssd1 vccd1 vccd1 _06962_/X sky130_fd_sc_hd__a21bo_1
XFILLER_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08701_ _08716_/A vssd1 vssd1 vccd1 vccd1 _08701_/X sky130_fd_sc_hd__clkbuf_2
X_09681_ _09684_/A vssd1 vssd1 vccd1 vccd1 _09886_/A sky130_fd_sc_hd__buf_1
X_06893_ _06893_/A vssd1 vssd1 vccd1 vccd1 _13187_/D sky130_fd_sc_hd__inv_2
XFILLER_67_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08632_ _08638_/A vssd1 vssd1 vccd1 vccd1 _08632_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08563_ _08811_/A vssd1 vssd1 vccd1 vccd1 _08817_/A sky130_fd_sc_hd__inv_2
XPHY_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07514_ _07609_/A _07514_/B vssd1 vssd1 vccd1 vccd1 _13005_/D sky130_fd_sc_hd__nor2_1
XFILLER_74_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08494_ _08457_/X _08474_/X _08494_/C _08494_/D vssd1 vssd1 vccd1 vccd1 _08494_/X
+ sky130_fd_sc_hd__and4bb_2
XPHY_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07445_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07445_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07376_ _11428_/X _07368_/X _13052_/Q _07369_/X vssd1 vssd1 vccd1 vccd1 _13052_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09115_ _09115_/A vssd1 vssd1 vccd1 vccd1 _09115_/X sky130_fd_sc_hd__clkbuf_2
X_06327_ _06327_/A vssd1 vssd1 vccd1 vccd1 _06327_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_176_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09046_ _09051_/A _12159_/X vssd1 vssd1 vccd1 vccd1 _12570_/D sky130_fd_sc_hd__nor2b_1
X_06258_ _13272_/Q vssd1 vssd1 vccd1 vccd1 _06258_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06189_ _06169_/Y _06022_/X _06163_/X _06188_/X vssd1 vssd1 vccd1 vccd1 _13285_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09948_ _08780_/Y _09943_/X _06243_/X _09938_/X _09941_/X vssd1 vssd1 vccd1 vccd1
+ _09948_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_161_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09879_ _09879_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09880_/B sky130_fd_sc_hd__or2_1
XFILLER_79_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11910_ _12441_/Q _10656_/Y _12091_/S vssd1 vssd1 vccd1 vccd1 _11910_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _12890_/CLK _12890_/D _07982_/X vssd1 vssd1 vccd1 vccd1 _12890_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _09951_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _09183_/A _11771_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11772_/X sky130_fd_sc_hd__mux2_1
XPHY_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _13244_/Q _06425_/A _11041_/A _10717_/X _06430_/X vssd1 vssd1 vccd1 vccd1
+ _10782_/A sky130_fd_sc_hd__o221a_1
XPHY_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10654_ _12620_/Q _11909_/S vssd1 vssd1 vccd1 vccd1 _12143_/S sky130_fd_sc_hd__nand2_8
XFILLER_55_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10585_ _10585_/A vssd1 vssd1 vccd1 vccd1 _10586_/B sky130_fd_sc_hd__inv_2
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12324_ _12999_/CLK _12324_/D vssd1 vssd1 vccd1 vccd1 _12324_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_1_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12166_/A0
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12255_ _12782_/Q _12855_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12255_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11206_ vssd1 vssd1 vccd1 vccd1 _11206_/HI _11206_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12186_ _11036_/A _10702_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12186_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11137_ _10755_/A _11100_/X _13250_/Q _11107_/X _11108_/X vssd1 vssd1 vccd1 vccd1
+ _11137_/X sky130_fd_sc_hd__a221o_2
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11068_ _10699_/X _10750_/X _06400_/X _10751_/X _10752_/X vssd1 vssd1 vccd1 vccd1
+ _11068_/X sky130_fd_sc_hd__a221o_1
XFILLER_95_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10019_ _12877_/Q vssd1 vssd1 vccd1 vccd1 _10019_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07230_ _07236_/A vssd1 vssd1 vccd1 vccd1 _07230_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07161_ _07161_/A vssd1 vssd1 vccd1 vccd1 _07161_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_145_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06112_ _12721_/Q vssd1 vssd1 vccd1 vccd1 _06112_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07092_ _09984_/A _09986_/B _09302_/A vssd1 vssd1 vccd1 vccd1 _10090_/A sky130_fd_sc_hd__or3_4
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput501 _11250_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput512 _11260_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__clkbuf_2
X_06043_ _12741_/Q _12709_/Q _06041_/Y _06042_/Y vssd1 vssd1 vccd1 vccd1 _06045_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput523 _11270_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__clkbuf_2
Xoutput534 _11280_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__clkbuf_2
Xoutput545 _11290_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__clkbuf_2
Xoutput556 _11300_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput567 _11310_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__clkbuf_2
Xoutput578 _12295_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_141_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput589 _12561_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__clkbuf_2
X_09802_ _09802_/A _09802_/B vssd1 vssd1 vccd1 vccd1 _09824_/A sky130_fd_sc_hd__or2_1
XFILLER_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07994_ _12887_/Q _07974_/X _07993_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _12887_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ _09733_/A vssd1 vssd1 vccd1 vccd1 _09733_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06945_ _12055_/X _06944_/Y _12055_/X _06944_/Y vssd1 vssd1 vccd1 vccd1 _06945_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_86_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09664_ _13199_/Q _13198_/Q _06792_/Y _06796_/Y vssd1 vssd1 vccd1 vccd1 _09666_/A
+ sky130_fd_sc_hd__o22a_1
X_06876_ _06874_/X _06875_/X _06874_/X _06875_/X vssd1 vssd1 vccd1 vccd1 _06876_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08615_ _08623_/A vssd1 vssd1 vccd1 vccd1 _08615_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09595_ _13157_/Q vssd1 vssd1 vccd1 vccd1 _09595_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_71_wb_clk_i _12960_/CLK vssd1 vssd1 vccd1 vccd1 _12955_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08546_ _12752_/Q vssd1 vssd1 vccd1 vccd1 _08546_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08477_ _13071_/Q _10395_/A _13066_/Q _07868_/Y vssd1 vssd1 vccd1 vccd1 _08482_/B
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07428_ _07428_/A vssd1 vssd1 vccd1 vccd1 _07428_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07359_ _11435_/X _07353_/X _13059_/Q _07354_/X vssd1 vssd1 vccd1 vccd1 _13059_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10370_ _10367_/B _10363_/A _10367_/A vssd1 vssd1 vccd1 vccd1 _10371_/C sky130_fd_sc_hd__o21a_1
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09029_ _09269_/A _09029_/B vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__or2_1
XFILLER_191_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12040_ _10783_/X _10784_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _12040_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12942_ _12942_/CLK _12942_/D _07744_/X vssd1 vssd1 vccd1 vccd1 _12942_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _12892_/CLK _12873_/D _08032_/X vssd1 vssd1 vccd1 vccd1 _12873_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11824_ _09905_/Y _12849_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11824_/X sky130_fd_sc_hd__mux2_1
XPHY_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11755_ _12100_/X _12473_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11755_/X sky130_fd_sc_hd__mux2_1
XPHY_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10706_ _13239_/Q _11083_/A _10686_/X _06982_/A _06537_/Y vssd1 vssd1 vccd1 vccd1
+ _11049_/A sky130_fd_sc_hd__o221a_1
XPHY_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11686_ _11685_/X _11404_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12385_/D sky130_fd_sc_hd__mux2_1
XPHY_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10637_ _08927_/A _08927_/B _10636_/Y vssd1 vssd1 vccd1 vccd1 _10637_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10568_ _10521_/A _09411_/Y _09423_/Y _10567_/Y _11390_/S vssd1 vssd1 vccd1 vccd1
+ _10568_/X sky130_fd_sc_hd__o311a_1
XFILLER_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12307_ _12975_/CLK _12307_/D vssd1 vssd1 vccd1 vccd1 _12307_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10499_ _12504_/Q _09143_/B _09144_/B vssd1 vssd1 vccd1 vccd1 _10499_/X sky130_fd_sc_hd__a21bo_1
XFILLER_154_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12238_ _12237_/X _12639_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12238_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ _12169_/A0 _08274_/X _13075_/Q vssd1 vssd1 vccd1 vccd1 _12169_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_1
X_06730_ _12009_/X _12035_/X _06724_/X _06725_/X _06729_/X vssd1 vssd1 vccd1 vccd1
+ _06730_/X sky130_fd_sc_hd__o32a_2
XFILLER_7_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06661_ _06658_/X _06659_/Y _06608_/X _06660_/X vssd1 vssd1 vccd1 vccd1 _13213_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08400_ _08402_/A vssd1 vssd1 vccd1 vccd1 _08417_/A sky130_fd_sc_hd__buf_2
X_09380_ _09379_/Y _12408_/Q _09336_/Y _12404_/Q vssd1 vssd1 vccd1 vccd1 _09380_/X
+ sky130_fd_sc_hd__o22a_1
X_06592_ _06589_/X _06590_/X _12171_/X _06591_/X vssd1 vssd1 vccd1 vccd1 _06592_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_33_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08331_ _12814_/Q _11589_/X _08335_/S vssd1 vssd1 vccd1 vccd1 _12814_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08262_ _08282_/A vssd1 vssd1 vccd1 vccd1 _08262_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07213_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07213_/X sky130_fd_sc_hd__clkbuf_1
X_08193_ _13112_/Q vssd1 vssd1 vccd1 vccd1 _08193_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07144_ _07152_/A vssd1 vssd1 vccd1 vccd1 _07144_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07075_ _07069_/X _07074_/X _06336_/Y _13150_/Q _07042_/A vssd1 vssd1 vccd1 vccd1
+ _13150_/D sky130_fd_sc_hd__a32o_1
XFILLER_69_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06026_ _12745_/Q vssd1 vssd1 vccd1 vccd1 _06026_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput375 _11161_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__clkbuf_2
Xoutput386 _11171_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput397 _11181_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07977_ _07998_/A vssd1 vssd1 vccd1 vccd1 _07977_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09716_ _09674_/Y _09748_/A _09715_/Y vssd1 vssd1 vccd1 vccd1 _09717_/B sky130_fd_sc_hd__o21a_1
X_06928_ _06926_/X _06927_/X _06926_/X _06927_/X vssd1 vssd1 vccd1 vccd1 _06928_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_43_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09647_ _09952_/A _09949_/A _09714_/C _09646_/B _09659_/B vssd1 vssd1 vccd1 vccd1
+ _09647_/X sky130_fd_sc_hd__a221o_2
XFILLER_71_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06859_ _06863_/A vssd1 vssd1 vccd1 vccd1 _06859_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09578_ _09578_/A _09578_/B _09578_/C vssd1 vssd1 vccd1 vccd1 _09592_/A sky130_fd_sc_hd__nor3_4
XFILLER_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08519_/X _12240_/X _06396_/A _12757_/Q vssd1 vssd1 vccd1 vccd1 _12757_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ _12829_/Q _10792_/A _11543_/S vssd1 vssd1 vccd1 vccd1 _11540_/X sky130_fd_sc_hd__mux2_1
XPHY_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ _12914_/Q _09180_/A _11481_/S vssd1 vssd1 vccd1 vccd1 _11471_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13210_ _13213_/CLK _13210_/D _06685_/X vssd1 vssd1 vccd1 vccd1 _13210_/Q sky130_fd_sc_hd__dfrtp_1
X_10422_ _12811_/Q _10422_/B vssd1 vssd1 vccd1 vccd1 _10429_/C sky130_fd_sc_hd__nand2_2
XFILLER_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10353_ _10357_/C vssd1 vssd1 vccd1 vccd1 _10355_/B sky130_fd_sc_hd__inv_2
X_13141_ _12168_/X _13141_/D _07125_/X vssd1 vssd1 vccd1 vccd1 _13141_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ _12165_/X _13072_/D _07326_/X vssd1 vssd1 vccd1 vccd1 _13072_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10284_ _12890_/Q vssd1 vssd1 vccd1 vccd1 _10284_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12023_ _11119_/X _11109_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _12023_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12925_ _13004_/CLK _12925_/D vssd1 vssd1 vccd1 vccd1 _12925_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _13257_/CLK _12856_/D _08077_/X vssd1 vssd1 vccd1 vccd1 _12856_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_73_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11806_/X _12071_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12445_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _12871_/CLK _12787_/D _08397_/X vssd1 vssd1 vccd1 vccd1 _12787_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11738_ _11737_/X _11367_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12444_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11669_ _11392_/X _09186_/A _11675_/S vssd1 vssd1 vccd1 vccd1 _11669_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07900_ _12921_/Q _11510_/X _07904_/S vssd1 vssd1 vccd1 vccd1 _12921_/D sky130_fd_sc_hd__mux2_1
XFILLER_102_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08880_ _08882_/A vssd1 vssd1 vccd1 vccd1 _08880_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07831_ _07827_/Y _12910_/Q _13026_/Q _10368_/A _07830_/X vssd1 vssd1 vccd1 vccd1
+ _07842_/B sky130_fd_sc_hd__a221o_1
XFILLER_97_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07762_ _12588_/Q _07762_/B vssd1 vssd1 vccd1 vccd1 _07763_/B sky130_fd_sc_hd__or2_1
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09501_ _09500_/A _09500_/B _09500_/Y vssd1 vssd1 vccd1 vccd1 _09502_/B sky130_fd_sc_hd__a21oi_1
X_06713_ _06672_/Y _12051_/X _06672_/Y _12051_/X vssd1 vssd1 vccd1 vccd1 _06720_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_07693_ _07705_/A vssd1 vssd1 vccd1 vccd1 _07693_/X sky130_fd_sc_hd__buf_2
XFILLER_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09432_ _09353_/X _09371_/X _09382_/X _09402_/Y _09431_/X vssd1 vssd1 vccd1 vccd1
+ _12450_/D sky130_fd_sc_hd__a311oi_4
X_06644_ _06641_/X _06642_/X _11897_/X _06643_/X vssd1 vssd1 vccd1 vccd1 _06644_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_92_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09363_ _12545_/Q vssd1 vssd1 vccd1 vccd1 _09363_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06575_ _06580_/A vssd1 vssd1 vccd1 vccd1 _06575_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08314_ _08325_/A vssd1 vssd1 vccd1 vccd1 _08314_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09294_ _10527_/A _10527_/B _09434_/B _09294_/D vssd1 vssd1 vccd1 vccd1 _09296_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_123_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08245_ _08199_/Y _08117_/X _13113_/Q _08122_/Y _08244_/Y vssd1 vssd1 vccd1 vccd1
+ _08246_/D sky130_fd_sc_hd__o221a_1
XFILLER_192_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08176_ _12804_/Q vssd1 vssd1 vccd1 vccd1 _08176_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07127_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07127_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07058_ _07074_/A vssd1 vssd1 vccd1 vccd1 _07058_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06009_ _09043_/A _09043_/B _11967_/S vssd1 vssd1 vccd1 vccd1 _06011_/A sky130_fd_sc_hd__or3_1
XFILLER_121_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10971_ _10969_/Y _10970_/Y _12537_/Q _12349_/Q vssd1 vssd1 vccd1 vccd1 _10976_/B
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_opt_3_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12710_ _12713_/CLK _12710_/D _08678_/X vssd1 vssd1 vccd1 vccd1 _12710_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12641_ _12870_/CLK _12641_/D _08866_/X vssd1 vssd1 vccd1 vccd1 _12641_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ _12977_/CLK _12572_/D vssd1 vssd1 vccd1 vccd1 _12572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11523_ _12812_/Q _09183_/A _11533_/S vssd1 vssd1 vccd1 vccd1 _11523_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11454_ _12897_/Q _09186_/A _11459_/S vssd1 vssd1 vccd1 vccd1 _11454_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ _10405_/A vssd1 vssd1 vccd1 vccd1 _10405_/Y sky130_fd_sc_hd__inv_2
X_11385_ _10583_/Y _12402_/D _11392_/S vssd1 vssd1 vccd1 vccd1 _11385_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13124_ _12168_/X _13124_/D _07167_/X vssd1 vssd1 vccd1 vccd1 _13124_/Q sky130_fd_sc_hd__dfrtp_2
X_10336_ _07804_/X _10335_/B _10342_/C _10320_/X vssd1 vssd1 vccd1 vccd1 _10336_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13055_ _12165_/X _13055_/D _07367_/X vssd1 vssd1 vccd1 vccd1 _13055_/Q sky130_fd_sc_hd__dfrtp_4
X_10267_ _12873_/Q vssd1 vssd1 vccd1 vccd1 _10267_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12006_ _11109_/X _11101_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10198_ _12780_/Q vssd1 vssd1 vccd1 vccd1 _10198_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12908_ _12166_/X _12908_/D _07929_/X vssd1 vssd1 vccd1 vccd1 _12908_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_128_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13269_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12839_ _12169_/A0 _12839_/D _08260_/X vssd1 vssd1 vccd1 vccd1 _12839_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06360_ _06370_/A vssd1 vssd1 vccd1 vccd1 _06360_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06291_ _06291_/A vssd1 vssd1 vccd1 vccd1 _06291_/Y sky130_fd_sc_hd__clkinv_4
X_08030_ _08036_/A vssd1 vssd1 vccd1 vccd1 _08030_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput30 io_in[36] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_1
Xinput41 la_data_in[101] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_1
Xinput52 la_data_in[111] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_1
Xinput63 la_data_in[121] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_1
XFILLER_162_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput74 la_data_in[16] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_1
Xinput85 la_data_in[26] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__buf_1
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
Xinput96 la_data_in[36] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__buf_1
XFILLER_196_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09981_ _09981_/A _09982_/D _09981_/C vssd1 vssd1 vccd1 vccd1 _10163_/A sky130_fd_sc_hd__or3_4
XFILLER_170_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08932_ _12424_/Q _08932_/B _12321_/Q vssd1 vssd1 vccd1 vccd1 _12620_/D sky130_fd_sc_hd__and3_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08863_ _08849_/X _06327_/Y _08852_/X _12643_/Q vssd1 vssd1 vccd1 vccd1 _12643_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater620 _11459_/S vssd1 vssd1 vccd1 vccd1 _11469_/S sky130_fd_sc_hd__buf_4
X_07814_ _13030_/Q vssd1 vssd1 vccd1 vccd1 _07814_/Y sky130_fd_sc_hd__inv_2
Xrepeater631 _11981_/S vssd1 vssd1 vccd1 vccd1 _12159_/S sky130_fd_sc_hd__buf_8
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater642 input339/X vssd1 vssd1 vccd1 vccd1 _09180_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_84_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08794_ _12670_/Q vssd1 vssd1 vccd1 vccd1 _08794_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07745_ _12615_/Q vssd1 vssd1 vccd1 vccd1 _08849_/A sky130_fd_sc_hd__inv_2
XFILLER_53_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07676_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07676_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09415_ _12402_/D vssd1 vssd1 vccd1 vccd1 _09415_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06627_ _06526_/X _06620_/B _06625_/Y _06556_/X _06626_/Y vssd1 vssd1 vccd1 vccd1
+ _06628_/A sky130_fd_sc_hd__o32a_1
XFILLER_52_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _12411_/Q vssd1 vssd1 vccd1 vccd1 _09346_/Y sky130_fd_sc_hd__inv_2
X_06558_ _06526_/X _06552_/B _06555_/Y _06556_/X _09798_/A vssd1 vssd1 vccd1 vccd1
+ _06559_/A sky130_fd_sc_hd__o32a_1
XFILLER_194_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09277_ _09283_/B _09277_/B _09277_/C _09286_/A vssd1 vssd1 vccd1 vccd1 _09278_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06489_ _06769_/A vssd1 vssd1 vccd1 vccd1 _06489_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08228_ _13097_/Q _10444_/A _13110_/Q _10480_/A vssd1 vssd1 vccd1 vccd1 _08232_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08159_ _13122_/Q vssd1 vssd1 vccd1 vccd1 _08159_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11170_ vssd1 vssd1 vccd1 vccd1 _11170_/HI _11170_/LO sky130_fd_sc_hd__conb_1
XFILLER_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10121_ _12849_/Q vssd1 vssd1 vccd1 vccd1 _10121_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10052_ _10052_/A _10796_/A vssd1 vssd1 vccd1 vccd1 _10052_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10954_ _10952_/Y _10953_/Y _12534_/Q _12346_/Q vssd1 vssd1 vccd1 vccd1 _10977_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10885_ _12525_/Q _12337_/Q _10884_/Y vssd1 vssd1 vccd1 vccd1 _10888_/D sky130_fd_sc_hd__a21o_1
XFILLER_32_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12624_ _12765_/CLK _12624_/D _08910_/X vssd1 vssd1 vccd1 vccd1 _12624_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12555_ _12558_/CLK _12555_/D vssd1 vssd1 vccd1 vccd1 _12555_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ _10384_/X _10792_/B _11513_/S vssd1 vssd1 vccd1 vccd1 _11506_/X sky130_fd_sc_hd__mux2_1
XPHY_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12486_ _12490_/CLK _12486_/D vssd1 vssd1 vccd1 vccd1 _12486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11437_ _12912_/Q _09180_/C _11443_/S vssd1 vssd1 vccd1 vccd1 _11437_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ _10661_/Y _12425_/Q _12103_/S vssd1 vssd1 vccd1 vccd1 _11368_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13107_ _12167_/X _13107_/D _07217_/X vssd1 vssd1 vccd1 vccd1 _13107_/Q sky130_fd_sc_hd__dfrtp_1
X_10319_ _10324_/A vssd1 vssd1 vccd1 vccd1 _10372_/A sky130_fd_sc_hd__inv_2
XFILLER_112_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11299_ vssd1 vssd1 vccd1 vccd1 _11299_/HI _11299_/LO sky130_fd_sc_hd__conb_1
XFILLER_140_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13038_ _12164_/X _13038_/D _07420_/X vssd1 vssd1 vccd1 vccd1 _13038_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07530_ _07532_/A vssd1 vssd1 vccd1 vccd1 _07531_/A sky130_fd_sc_hd__inv_2
XFILLER_19_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07461_ _11463_/X _07459_/X _13022_/Q _07460_/X vssd1 vssd1 vccd1 vccd1 _13022_/D
+ sky130_fd_sc_hd__a22o_1
X_09200_ _09216_/A vssd1 vssd1 vccd1 vccd1 _09200_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06412_ _06412_/A vssd1 vssd1 vccd1 vccd1 _06412_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07392_ _11422_/X _07384_/X _13046_/Q _07385_/X vssd1 vssd1 vccd1 vccd1 _13046_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06343_ _07742_/B _06314_/X _06342_/Y _13257_/Q _06306_/A vssd1 vssd1 vccd1 vccd1
+ _13257_/D sky130_fd_sc_hd__a32o_1
X_09131_ _12511_/Q _09115_/A _07566_/X _09116_/A vssd1 vssd1 vccd1 vccd1 _12511_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09062_ _10227_/A _12145_/X vssd1 vssd1 vccd1 vccd1 _12556_/D sky130_fd_sc_hd__nor2b_4
XFILLER_33_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06274_ _06269_/X _06247_/X _06271_/Y _13270_/Q _06273_/X vssd1 vssd1 vccd1 vccd1
+ _13270_/D sky130_fd_sc_hd__a32o_1
XFILLER_120_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_96_wb_clk_i _13235_/CLK vssd1 vssd1 vccd1 vccd1 _13177_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08013_ _12880_/Q _07996_/A _07300_/X _07998_/A vssd1 vssd1 vccd1 vccd1 _12880_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12441_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09964_ _09981_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _11981_/S sky130_fd_sc_hd__nor2_8
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08915_ _08962_/A vssd1 vssd1 vccd1 vccd1 _08915_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09895_ _09890_/Y _07732_/X _06346_/A _09892_/X _09894_/X vssd1 vssd1 vccd1 vccd1
+ _09895_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08846_ _08851_/A vssd1 vssd1 vccd1 vccd1 _08846_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08777_ _12675_/Q vssd1 vssd1 vccd1 vccd1 _08777_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07728_ _07749_/A vssd1 vssd1 vccd1 vccd1 _07728_/X sky130_fd_sc_hd__clkbuf_1
XPHY_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07659_ _07659_/A _12961_/Q vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__nand2_1
XPHY_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10670_ _12433_/Q vssd1 vssd1 vccd1 vccd1 _10670_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09329_ _09329_/A _09329_/B vssd1 vssd1 vccd1 vccd1 _10541_/A sky130_fd_sc_hd__or2_1
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12340_ _12357_/CLK _12340_/D vssd1 vssd1 vccd1 vccd1 _12340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12271_ _10133_/X _12897_/Q _11863_/X _11864_/X _11348_/X _11348_/S vssd1 vssd1 vccd1
+ vccd1 _12287_/D sky130_fd_sc_hd__mux4_2
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11222_ vssd1 vssd1 vccd1 vccd1 _11222_/HI _11222_/LO sky130_fd_sc_hd__conb_1
XFILLER_175_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11153_ vssd1 vssd1 vccd1 vccd1 _11153_/HI _11153_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10104_ _12775_/Q vssd1 vssd1 vccd1 vccd1 _10104_/Y sky130_fd_sc_hd__inv_2
X_11084_ _12089_/X vssd1 vssd1 vccd1 vccd1 _11084_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput220 la_oenb[32] vssd1 vssd1 vccd1 vccd1 input220/X sky130_fd_sc_hd__buf_1
XFILLER_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput231 la_oenb[42] vssd1 vssd1 vccd1 vccd1 input231/X sky130_fd_sc_hd__buf_1
Xinput242 la_oenb[52] vssd1 vssd1 vccd1 vccd1 input242/X sky130_fd_sc_hd__buf_1
XFILLER_48_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10035_ _10035_/A vssd1 vssd1 vccd1 vccd1 _10151_/A sky130_fd_sc_hd__clkbuf_4
Xinput253 la_oenb[62] vssd1 vssd1 vccd1 vccd1 input253/X sky130_fd_sc_hd__buf_1
XFILLER_49_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput264 la_oenb[72] vssd1 vssd1 vccd1 vccd1 input264/X sky130_fd_sc_hd__buf_1
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput275 la_oenb[82] vssd1 vssd1 vccd1 vccd1 input275/X sky130_fd_sc_hd__buf_1
Xinput286 la_oenb[92] vssd1 vssd1 vccd1 vccd1 input286/X sky130_fd_sc_hd__buf_1
XFILLER_84_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput297 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 input297/X sky130_fd_sc_hd__buf_1
XFILLER_1_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11986_ _11122_/X _11115_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _11986_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10937_ _12344_/Q vssd1 vssd1 vccd1 vccd1 _10937_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10868_ _10854_/Y _10855_/Y _10865_/X _10867_/Y vssd1 vssd1 vccd1 vccd1 _10890_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12607_ _13260_/CLK _12607_/D _08972_/X vssd1 vssd1 vccd1 vccd1 _12607_/Q sky130_fd_sc_hd__dfstp_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _10799_/A _10799_/B vssd1 vssd1 vccd1 vccd1 _10799_/Y sky130_fd_sc_hd__nor2_2
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12538_ _12540_/CLK _12538_/D vssd1 vssd1 vccd1 vccd1 _12538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12469_ _12472_/CLK _12469_/D vssd1 vssd1 vccd1 vccd1 _12469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06961_ _06961_/A _06961_/B vssd1 vssd1 vccd1 vccd1 _06961_/Y sky130_fd_sc_hd__nand2_1
X_08700_ _08715_/A vssd1 vssd1 vccd1 vccd1 _08700_/X sky130_fd_sc_hd__clkbuf_2
X_09680_ _09679_/Y _12613_/Q _12876_/Q _12614_/Q vssd1 vssd1 vccd1 vccd1 _09684_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_95_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06892_ _06841_/A _06883_/B _06890_/Y _06556_/X _06891_/Y vssd1 vssd1 vccd1 vccd1
+ _06893_/A sky130_fd_sc_hd__o32a_1
XFILLER_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_143_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12892_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08631_ _11938_/X _08624_/X _12729_/Q _08625_/X vssd1 vssd1 vccd1 vccd1 _12729_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ _11961_/X _08562_/B vssd1 vssd1 vccd1 vccd1 _08811_/A sky130_fd_sc_hd__or2_2
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07513_ _09227_/A _07497_/Y _07522_/B _11982_/X _07512_/Y vssd1 vssd1 vccd1 vccd1
+ _07514_/B sky130_fd_sc_hd__o32a_1
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08493_ _08484_/X _08493_/B _08493_/C _08493_/D vssd1 vssd1 vccd1 vccd1 _08494_/D
+ sky130_fd_sc_hd__and4b_1
XPHY_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07444_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07444_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07375_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07375_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09114_ _12524_/Q _09107_/X _07980_/X _09108_/X vssd1 vssd1 vccd1 vccd1 _12524_/D
+ sky130_fd_sc_hd__a22o_1
X_06326_ _06108_/B _06320_/Y _06108_/B _06320_/Y vssd1 vssd1 vccd1 vccd1 _06327_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06257_ _06280_/A vssd1 vssd1 vccd1 vccd1 _06257_/X sky130_fd_sc_hd__clkbuf_1
X_09045_ _10244_/A vssd1 vssd1 vccd1 vccd1 _09051_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06188_ _06035_/A _06187_/X _06035_/A _06187_/X vssd1 vssd1 vccd1 vccd1 _06188_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_2_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09947_ _08784_/Y _09943_/X _06248_/X _09938_/X _09941_/X vssd1 vssd1 vccd1 vccd1
+ _09947_/Y sky130_fd_sc_hd__o221ai_1
X_09878_ _09492_/X _09876_/Y _09877_/X _09700_/A vssd1 vssd1 vccd1 vccd1 _09878_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08829_ _08814_/A _08817_/X _06336_/Y _12657_/Q _08567_/A vssd1 vssd1 vccd1 vccd1
+ _12657_/D sky130_fd_sc_hd__a32o_1
XFILLER_79_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _09948_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11840_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _12115_/X _12477_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__mux2_1
XPHY_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _13244_/Q vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__inv_2
XFILLER_0_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10653_ _11907_/X _10653_/B vssd1 vssd1 vccd1 vccd1 _10653_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10584_ _10608_/A _10608_/B _12372_/Q vssd1 vssd1 vccd1 vccd1 _11404_/S sky130_fd_sc_hd__or3b_4
XFILLER_70_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12323_ _12995_/CLK _12323_/D vssd1 vssd1 vccd1 vccd1 _12323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12254_ _12253_/X _12647_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12254_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11205_ vssd1 vssd1 vccd1 vccd1 _11205_/HI _11205_/LO sky130_fd_sc_hd__conb_1
XFILLER_134_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12185_ _10700_/X _10697_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _12185_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11136_ _10736_/A _10759_/A _13252_/Q _11086_/A _12195_/X vssd1 vssd1 vccd1 vccd1
+ _11136_/X sky130_fd_sc_hd__a221o_1
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11067_ _11041_/X _11054_/X _06392_/X _11055_/X _11060_/X vssd1 vssd1 vccd1 vccd1
+ _11067_/X sky130_fd_sc_hd__a221o_1
XFILLER_114_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10018_ _10165_/A vssd1 vssd1 vccd1 vccd1 _10018_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11969_ _09299_/Y _09297_/Y _11969_/S vssd1 vssd1 vccd1 vccd1 _11969_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07160_ _07160_/A vssd1 vssd1 vccd1 vccd1 _07160_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06111_ _12722_/Q _12690_/Q _12722_/Q _12690_/Q vssd1 vssd1 vccd1 vccd1 _06125_/A
+ sky130_fd_sc_hd__o2bb2ai_1
X_07091_ _09984_/B vssd1 vssd1 vccd1 vccd1 _09986_/B sky130_fd_sc_hd__buf_2
XFILLER_173_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput502 _11251_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__clkbuf_2
X_06042_ _12709_/Q vssd1 vssd1 vccd1 vccd1 _06042_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput513 _11261_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput524 _11271_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__clkbuf_2
Xoutput535 _11281_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput546 _11291_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__clkbuf_2
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput557 _11301_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput568 _11311_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__clkbuf_2
Xoutput579 _12296_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09801_ _09800_/A _09800_/B _09800_/Y vssd1 vssd1 vccd1 vccd1 _09823_/A sky130_fd_sc_hd__a21o_1
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07993_ _07993_/A vssd1 vssd1 vccd1 vccd1 _07993_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09732_ _09747_/A _09825_/A _09711_/Y vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__a21oi_2
XFILLER_80_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06944_ _12053_/X vssd1 vssd1 vccd1 vccd1 _06944_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09663_ _06822_/Y _06830_/Y _09652_/Y _09653_/Y vssd1 vssd1 vccd1 vccd1 _09668_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_94_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06875_ _11997_/X _11994_/X _11997_/X _11994_/X vssd1 vssd1 vccd1 vccd1 _06875_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08614_ _11945_/X _08608_/X _12736_/Q _08610_/X vssd1 vssd1 vccd1 vccd1 _12736_/D
+ sky130_fd_sc_hd__a22o_1
X_09594_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09594_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08545_ _08569_/A vssd1 vssd1 vccd1 vccd1 _08545_/X sky130_fd_sc_hd__clkbuf_1
XPHY_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08476_ _13066_/Q _07868_/Y _08475_/Y _12898_/Q vssd1 vssd1 vccd1 vccd1 _08476_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07427_ _11476_/X _07412_/X _13035_/Q _07415_/X vssd1 vssd1 vccd1 vccd1 _13035_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_40_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12977_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07358_ _07360_/A vssd1 vssd1 vccd1 vccd1 _07358_/X sky130_fd_sc_hd__clkbuf_1
X_06309_ _06099_/Y _06100_/Y _06129_/A _06103_/B vssd1 vssd1 vccd1 vccd1 _06309_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07289_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07289_/X sky130_fd_sc_hd__clkbuf_1
X_09028_ _12303_/Q vssd1 vssd1 vccd1 vccd1 _09029_/B sky130_fd_sc_hd__inv_2
XFILLER_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ _13257_/CLK _12941_/D _07749_/X vssd1 vssd1 vccd1 vccd1 _12941_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12872_ _12872_/CLK _12872_/D _08034_/X vssd1 vssd1 vccd1 vccd1 _12872_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _09902_/Y _12848_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11823_/X sky130_fd_sc_hd__mux2_2
XFILLER_73_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11754_ _11753_/X _11376_/X _11774_/S vssd1 vssd1 vccd1 vccd1 _12428_/D sky130_fd_sc_hd__mux2_1
XPHY_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10705_ _13240_/Q _11083_/A _10693_/A _11075_/A _06537_/Y vssd1 vssd1 vccd1 vccd1
+ _11062_/A sky130_fd_sc_hd__o221a_1
XPHY_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11685_ _11404_/X _09244_/A _11691_/S vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__mux2_1
XPHY_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10636_ _10636_/A vssd1 vssd1 vccd1 vccd1 _10636_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10567_ _10521_/A _09411_/Y _09423_/Y vssd1 vssd1 vccd1 vccd1 _10567_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ _12939_/CLK _12306_/D vssd1 vssd1 vccd1 vccd1 _12306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13286_ _13286_/CLK _13286_/D _11147_/X vssd1 vssd1 vccd1 vccd1 _13286_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10498_ _12503_/Q _09142_/B _09143_/B vssd1 vssd1 vccd1 vccd1 _10498_/X sky130_fd_sc_hd__a21bo_1
X_12237_ _12773_/Q _12846_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12168_ _12168_/A0 input32/X hold1/A vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11119_ _11041_/X _11100_/X _13244_/Q _11107_/X _11108_/X vssd1 vssd1 vccd1 vccd1
+ _11119_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12099_ _12098_/X _12429_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12099_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput6 io_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_1
XFILLER_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06660_ _06652_/X _06653_/X _06652_/X _06653_/X vssd1 vssd1 vccd1 vccd1 _06660_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06591_ _06589_/X _06590_/X _06589_/X _06590_/X vssd1 vssd1 vccd1 vccd1 _06591_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08330_ _08339_/A vssd1 vssd1 vccd1 vccd1 _08330_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_189_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08261_ _12839_/Q _08251_/X _07300_/X _11417_/S vssd1 vssd1 vccd1 vccd1 _12839_/D
+ sky130_fd_sc_hd__a22o_1
X_07212_ _11575_/X _07201_/X _13110_/Q _07204_/X vssd1 vssd1 vccd1 vccd1 _13110_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08192_ _09009_/A vssd1 vssd1 vccd1 vccd1 _09019_/A sky130_fd_sc_hd__buf_4
XFILLER_118_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07143_ _11535_/X _07130_/X _13134_/Q _07131_/X vssd1 vssd1 vccd1 vccd1 _13134_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07074_ _07074_/A vssd1 vssd1 vccd1 vccd1 _07074_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06025_ _06025_/A _06025_/B vssd1 vssd1 vccd1 vccd1 _06025_/X sky130_fd_sc_hd__or2_1
XFILLER_126_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput376 _11162_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__clkbuf_2
Xoutput387 _11172_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput398 _11155_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07976_ _07976_/A vssd1 vssd1 vccd1 vccd1 _07998_/A sky130_fd_sc_hd__inv_2
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09715_ _09669_/Y _09671_/Y _09694_/Y vssd1 vssd1 vccd1 vccd1 _09715_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06927_ _12001_/X _11998_/X _12001_/X _11998_/X vssd1 vssd1 vccd1 vccd1 _06927_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09646_ _09714_/C _09646_/B vssd1 vssd1 vccd1 vccd1 _09659_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06858_ _06829_/X _06844_/Y _06769_/X _06857_/Y vssd1 vssd1 vccd1 vccd1 _13192_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09577_ _09576_/A _09576_/B _09576_/Y vssd1 vssd1 vccd1 vccd1 _09578_/C sky130_fd_sc_hd__a21o_1
X_06789_ _06787_/X _06788_/X _06787_/X _06788_/X vssd1 vssd1 vccd1 vccd1 _06789_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _08533_/A vssd1 vssd1 vccd1 vccd1 _08528_/X sky130_fd_sc_hd__clkbuf_1
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ _13062_/Q _10373_/A _13057_/Q _10357_/A vssd1 vssd1 vccd1 vccd1 _08459_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11470_ _12913_/Q _09180_/B _11481_/S vssd1 vssd1 vccd1 vccd1 _11470_/X sky130_fd_sc_hd__mux2_1
XPHY_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10421_ _10420_/A _10420_/B _10422_/B _10411_/A vssd1 vssd1 vccd1 vccd1 _10421_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_137_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13140_ _12168_/X _13140_/D _07127_/X vssd1 vssd1 vccd1 vccd1 _13140_/Q sky130_fd_sc_hd__dfrtp_1
X_10352_ _10352_/A _10352_/B _10352_/C vssd1 vssd1 vccd1 vccd1 _10357_/C sky130_fd_sc_hd__or3_4
XFILLER_125_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _12165_/X _13071_/D _07328_/X vssd1 vssd1 vccd1 vccd1 _13071_/Q sky130_fd_sc_hd__dfrtp_4
X_10283_ _12785_/Q vssd1 vssd1 vccd1 vccd1 _10283_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12022_ _11098_/X _11093_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12022_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12924_ _12166_/X _12924_/D _07793_/X vssd1 vssd1 vccd1 vccd1 _12924_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12855_ _12890_/CLK _12855_/D _08079_/X vssd1 vssd1 vccd1 vccd1 _12855_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11806_ _12071_/X _11805_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11806_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12892_/CLK _12786_/D _08405_/X vssd1 vssd1 vccd1 vccd1 _12786_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11367_/X _11736_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11737_/X sky130_fd_sc_hd__mux2_1
XPHY_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11668_ _11667_/X _11379_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12376_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10619_ _10619_/A _10619_/B vssd1 vssd1 vccd1 vccd1 _10620_/A sky130_fd_sc_hd__or2_1
XPHY_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11599_ _10461_/X _09180_/B _11603_/S vssd1 vssd1 vccd1 vccd1 _11599_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13269_ _13269_/CLK _13269_/D _06275_/X vssd1 vssd1 vccd1 vccd1 _13269_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07830_ _13015_/Q _10333_/A _13023_/Q _10357_/B vssd1 vssd1 vccd1 vccd1 _07830_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07761_ _12587_/Q _07761_/B vssd1 vssd1 vccd1 vccd1 _07762_/B sky130_fd_sc_hd__or2_1
XFILLER_65_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09500_ _09500_/A _09500_/B vssd1 vssd1 vccd1 vccd1 _09500_/Y sky130_fd_sc_hd__nor2_2
X_06712_ _06694_/A _06694_/B _06694_/X vssd1 vssd1 vccd1 vccd1 _06712_/X sky130_fd_sc_hd__a21bo_1
XFILLER_38_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07692_ _07717_/A vssd1 vssd1 vccd1 vccd1 _07705_/A sky130_fd_sc_hd__inv_2
XFILLER_38_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09431_ _09431_/A _09431_/B _09427_/X _09430_/X vssd1 vssd1 vccd1 vccd1 _09431_/X
+ sky130_fd_sc_hd__or4bb_4
X_06643_ _06641_/X _06642_/X _06641_/X _06642_/X vssd1 vssd1 vccd1 vccd1 _06643_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09362_ _12462_/Q vssd1 vssd1 vccd1 vccd1 _09362_/Y sky130_fd_sc_hd__inv_2
X_06574_ _06507_/X _09798_/B _06489_/X _06573_/Y vssd1 vssd1 vccd1 vccd1 _13222_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_166_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08313_ _08372_/A vssd1 vssd1 vccd1 vccd1 _08325_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09293_ _09293_/A _09293_/B _09293_/C _09293_/D vssd1 vssd1 vccd1 vccd1 _09294_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08244_ _13098_/Q _10455_/B vssd1 vssd1 vccd1 vccd1 _08244_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08175_ _08166_/X _08175_/B _08175_/C _08175_/D vssd1 vssd1 vccd1 vccd1 _08191_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_192_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07126_ _11542_/X _07113_/X _13141_/Q _07116_/X vssd1 vssd1 vccd1 vccd1 _13141_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07057_ _07063_/A vssd1 vssd1 vccd1 vccd1 _07057_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06008_ _12550_/Q vssd1 vssd1 vccd1 vccd1 _09433_/A sky130_fd_sc_hd__inv_2
XFILLER_86_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07959_ _07961_/A vssd1 vssd1 vccd1 vccd1 _07959_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10970_ _12349_/Q vssd1 vssd1 vccd1 vccd1 _10970_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09629_ _12874_/Q vssd1 vssd1 vccd1 vccd1 _09629_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12640_ _12870_/CLK _12640_/D _08869_/X vssd1 vssd1 vccd1 vccd1 _12640_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12571_ _12993_/CLK _12571_/D vssd1 vssd1 vccd1 vccd1 _12571_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11522_ _12811_/Q _09185_/A _11522_/S vssd1 vssd1 vccd1 vccd1 _11522_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11453_ _12896_/Q _09186_/B _11459_/S vssd1 vssd1 vccd1 vccd1 _11453_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10404_ _12804_/Q _10458_/A vssd1 vssd1 vccd1 vccd1 _10404_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11384_ _10565_/Y _12395_/D _11392_/S vssd1 vssd1 vccd1 vccd1 _11384_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13123_ _12168_/X _13123_/D _07171_/X vssd1 vssd1 vccd1 vccd1 _13123_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_194_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10335_ _12900_/Q _10335_/B vssd1 vssd1 vccd1 vccd1 _10342_/C sky130_fd_sc_hd__nand2_4
XFILLER_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13054_ _12165_/X _13054_/D _07371_/X vssd1 vssd1 vccd1 vccd1 _13054_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10266_ _12784_/Q vssd1 vssd1 vccd1 vccd1 _10266_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12005_ _11064_/X _10759_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12005_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10197_ _10195_/Y _10000_/A _10196_/Y _10137_/X vssd1 vssd1 vccd1 vccd1 _10197_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12907_ _12166_/X _12907_/D _07931_/X vssd1 vssd1 vccd1 vccd1 _12907_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12838_ _12840_/CLK _12838_/D _08262_/X vssd1 vssd1 vccd1 vccd1 _12838_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12769_ _12769_/CLK _12769_/D _08498_/X vssd1 vssd1 vccd1 vccd1 _12769_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06290_ _06180_/A _06289_/X _06180_/A _06289_/X vssd1 vssd1 vccd1 vccd1 _06291_/A
+ sky130_fd_sc_hd__a2bb2o_2
Xinput20 io_in[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_1
Xinput31 io_in[37] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_1
XFILLER_174_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput42 la_data_in[102] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_1
Xinput53 la_data_in[112] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_1
Xinput64 la_data_in[122] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_1
XFILLER_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput75 la_data_in[17] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_1
XFILLER_116_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput86 la_data_in[27] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__buf_1
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput97 la_data_in[37] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__buf_1
XFILLER_116_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09980_ _12892_/Q vssd1 vssd1 vccd1 vccd1 _09980_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08931_ _08931_/A vssd1 vssd1 vccd1 vccd1 _08932_/B sky130_fd_sc_hd__inv_2
XFILLER_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08862_ _08866_/A vssd1 vssd1 vccd1 vccd1 _08862_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_112_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater610 _11803_/S vssd1 vssd1 vccd1 vccd1 _11819_/S sky130_fd_sc_hd__buf_8
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07813_ _12916_/Q vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__inv_2
Xrepeater621 _07409_/Y vssd1 vssd1 vccd1 vccd1 _11459_/S sky130_fd_sc_hd__buf_6
XFILLER_85_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08793_ _08807_/A vssd1 vssd1 vccd1 vccd1 _08793_/X sky130_fd_sc_hd__clkbuf_1
Xrepeater632 input360/X vssd1 vssd1 vccd1 vccd1 _09243_/D sky130_fd_sc_hd__buf_8
Xrepeater643 input338/X vssd1 vssd1 vccd1 vccd1 _09180_/D sky130_fd_sc_hd__buf_6
XFILLER_42_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07744_ _07749_/A vssd1 vssd1 vccd1 vccd1 _07744_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07675_ _09279_/B vssd1 vssd1 vccd1 vccd1 _09283_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09414_ _12460_/Q _09411_/Y _09354_/Y _12400_/D _09413_/X vssd1 vssd1 vccd1 vccd1
+ _09422_/B sky130_fd_sc_hd__a221o_1
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06626_ _13216_/Q vssd1 vssd1 vccd1 vccd1 _06626_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ _09341_/Y _12410_/Q _12466_/Q _09342_/Y _09344_/X vssd1 vssd1 vccd1 vccd1
+ _09353_/B sky130_fd_sc_hd__a221oi_2
X_06557_ _13223_/Q vssd1 vssd1 vccd1 vccd1 _09798_/A sky130_fd_sc_hd__inv_2
XFILLER_194_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09276_ _10015_/B _09276_/B _09276_/C vssd1 vssd1 vccd1 vccd1 _09286_/A sky130_fd_sc_hd__or3_1
XFILLER_166_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06488_ _13229_/Q vssd1 vssd1 vccd1 vccd1 _06488_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08227_ _13105_/Q _10467_/A _08226_/Y _12805_/Q vssd1 vssd1 vccd1 vccd1 _08232_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08158_ _13132_/Q _10454_/B _13125_/Q _10433_/A vssd1 vssd1 vccd1 vccd1 _08162_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07109_ _11969_/S _09984_/B _09302_/A vssd1 vssd1 vccd1 vccd1 _09978_/B sky130_fd_sc_hd__or3_4
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08089_ _12852_/Q _08082_/X _07290_/X _08083_/X vssd1 vssd1 vccd1 vccd1 _12852_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_161_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10120_ _09510_/Y _10023_/X _10119_/Y _10025_/X vssd1 vssd1 vccd1 vccd1 _10128_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_134_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10051_ _10277_/A vssd1 vssd1 vccd1 vccd1 _10051_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10953_ _12346_/Q vssd1 vssd1 vccd1 vccd1 _10953_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10884_ _12525_/Q _12337_/Q vssd1 vssd1 vccd1 vccd1 _10884_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12623_ _12646_/CLK _12623_/D _08912_/X vssd1 vssd1 vccd1 vccd1 _12623_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ _12169_/A0 _12554_/D _09064_/X vssd1 vssd1 vccd1 vccd1 _12554_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_196_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11505_ _10383_/Y _09179_/C _11513_/S vssd1 vssd1 vccd1 vccd1 _11505_/X sky130_fd_sc_hd__mux2_1
XPHY_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12485_ _12485_/CLK _12485_/D vssd1 vssd1 vccd1 vccd1 _12485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11436_ _12911_/Q _09180_/D _11443_/S vssd1 vssd1 vccd1 vccd1 _11436_/X sky130_fd_sc_hd__mux2_1
X_11367_ _11366_/X _12444_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _11367_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13106_ _12167_/X _13106_/D _07221_/X vssd1 vssd1 vccd1 vccd1 _13106_/Q sky130_fd_sc_hd__dfrtp_1
X_10318_ _10318_/A vssd1 vssd1 vccd1 vccd1 _10318_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11298_ vssd1 vssd1 vccd1 vccd1 _11298_/HI _11298_/LO sky130_fd_sc_hd__conb_1
XFILLER_112_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13037_ _12164_/X _13037_/D _07422_/X vssd1 vssd1 vccd1 vccd1 _13037_/Q sky130_fd_sc_hd__dfrtp_1
X_10249_ _12856_/Q vssd1 vssd1 vccd1 vccd1 _10249_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07460_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07460_/X sky130_fd_sc_hd__buf_2
XFILLER_50_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06411_ _06403_/X _12204_/X _06396_/X _06410_/X vssd1 vssd1 vccd1 vccd1 _13239_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07391_ _07391_/A vssd1 vssd1 vccd1 vccd1 _07391_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_188_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ _12512_/Q _09123_/X _07564_/X _09124_/X vssd1 vssd1 vccd1 vccd1 _12512_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06342_ _06342_/A vssd1 vssd1 vccd1 vccd1 _06342_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09061_ _10227_/A _12146_/X vssd1 vssd1 vccd1 vccd1 _12557_/D sky130_fd_sc_hd__nor2b_4
X_06273_ _06306_/A vssd1 vssd1 vccd1 vccd1 _06273_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08012_ _08018_/A vssd1 vssd1 vccd1 vccd1 _08012_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09963_ _11967_/S vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_65_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12937_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08914_ _08963_/A vssd1 vssd1 vccd1 vccd1 _08962_/A sky130_fd_sc_hd__clkbuf_4
X_09894_ _12878_/Q _09910_/B vssd1 vssd1 vccd1 vccd1 _09894_/X sky130_fd_sc_hd__or2_1
XFILLER_98_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08845_ _07746_/X _06291_/Y _08837_/X _12650_/Q vssd1 vssd1 vccd1 vccd1 _12650_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08776_ _08789_/A vssd1 vssd1 vccd1 vccd1 _08776_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07727_ _12946_/Q _07717_/X _07698_/X _07726_/Y _09288_/A vssd1 vssd1 vccd1 vccd1
+ _12946_/D sky130_fd_sc_hd__o221a_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07658_ _07658_/A _07658_/B _07658_/C vssd1 vssd1 vccd1 vccd1 _07668_/B sky130_fd_sc_hd__nor3_4
XPHY_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06609_ _11893_/X _11898_/X vssd1 vssd1 vccd1 vccd1 _06609_/X sky130_fd_sc_hd__or2_1
XFILLER_198_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07589_ _12301_/Q vssd1 vssd1 vccd1 vccd1 _09284_/B sky130_fd_sc_hd__inv_2
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09328_ _09328_/A _09328_/B vssd1 vssd1 vccd1 vccd1 _09329_/B sky130_fd_sc_hd__or2_1
XFILLER_185_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09259_ _09259_/A vssd1 vssd1 vccd1 vccd1 _09259_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _10115_/Y _12896_/Q _11861_/X _11862_/X _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12286_/D sky130_fd_sc_hd__mux4_2
XFILLER_181_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11221_ vssd1 vssd1 vccd1 vccd1 _11221_/HI _11221_/LO sky130_fd_sc_hd__conb_1
XFILLER_153_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11152_ vssd1 vssd1 vccd1 vccd1 _11152_/HI _11152_/LO sky130_fd_sc_hd__conb_1
XFILLER_175_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10103_ _13258_/Q vssd1 vssd1 vccd1 vccd1 _10103_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11083_ _11083_/A vssd1 vssd1 vccd1 vccd1 _11083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput210 la_oenb[23] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__buf_1
XFILLER_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput221 la_oenb[33] vssd1 vssd1 vccd1 vccd1 input221/X sky130_fd_sc_hd__buf_1
Xinput232 la_oenb[43] vssd1 vssd1 vccd1 vccd1 input232/X sky130_fd_sc_hd__buf_1
XFILLER_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10034_ _10034_/A vssd1 vssd1 vccd1 vccd1 _10792_/D sky130_fd_sc_hd__buf_2
XFILLER_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput243 la_oenb[53] vssd1 vssd1 vccd1 vccd1 input243/X sky130_fd_sc_hd__buf_1
XFILLER_0_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput254 la_oenb[63] vssd1 vssd1 vccd1 vccd1 input254/X sky130_fd_sc_hd__buf_1
Xinput265 la_oenb[73] vssd1 vssd1 vccd1 vccd1 input265/X sky130_fd_sc_hd__buf_1
XFILLER_76_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput276 la_oenb[83] vssd1 vssd1 vccd1 vccd1 input276/X sky130_fd_sc_hd__buf_1
Xinput287 la_oenb[93] vssd1 vssd1 vccd1 vccd1 input287/X sky130_fd_sc_hd__buf_1
XFILLER_29_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput298 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 input298/X sky130_fd_sc_hd__buf_1
XFILLER_64_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11985_ _11126_/X _11119_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _11985_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10936_ _12532_/Q vssd1 vssd1 vccd1 vccd1 _10936_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10867_ _12519_/Q _12331_/Q _10866_/X _10851_/X _10858_/A vssd1 vssd1 vccd1 vccd1
+ _10867_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_32_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12606_ _13244_/CLK _12606_/D vssd1 vssd1 vccd1 vccd1 _12606_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _12322_/Q vssd1 vssd1 vccd1 vccd1 _10799_/B sky130_fd_sc_hd__inv_2
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12537_ _12537_/CLK _12537_/D vssd1 vssd1 vccd1 vccd1 _12537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12468_ _12468_/CLK _12468_/D vssd1 vssd1 vccd1 vccd1 _12468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11419_ _12894_/Q _09185_/D _11449_/S vssd1 vssd1 vccd1 vccd1 _11419_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12399_ _12985_/CLK _12399_/D vssd1 vssd1 vccd1 vccd1 _12399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06960_ _11854_/X _06960_/B vssd1 vssd1 vccd1 vccd1 _06961_/B sky130_fd_sc_hd__or2_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06891_ _13187_/Q vssd1 vssd1 vccd1 vccd1 _06891_/Y sky130_fd_sc_hd__inv_2
X_08630_ _08638_/A vssd1 vssd1 vccd1 vccd1 _08630_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08561_ _12750_/Q vssd1 vssd1 vccd1 vccd1 _08561_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07512_ _13005_/Q vssd1 vssd1 vccd1 vccd1 _07512_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08492_ _13042_/Q _07822_/Y _13062_/Q _10373_/A _08491_/X vssd1 vssd1 vccd1 vccd1
+ _08493_/D sky130_fd_sc_hd__o221a_1
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_112_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 _12747_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07443_ _07443_/A vssd1 vssd1 vccd1 vccd1 _07443_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07374_ _11429_/X _07368_/X _13053_/Q _07369_/X vssd1 vssd1 vccd1 vccd1 _13053_/D
+ sky130_fd_sc_hd__a22o_1
X_09113_ _12525_/Q _09107_/X _07975_/X _09108_/X vssd1 vssd1 vccd1 vccd1 _12525_/D
+ sky130_fd_sc_hd__a22o_1
X_06325_ _06344_/A vssd1 vssd1 vccd1 vccd1 _06325_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09044_ _12312_/Q _10190_/A vssd1 vssd1 vccd1 vccd1 _10244_/A sky130_fd_sc_hd__or2_4
XFILLER_135_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06256_ _06252_/Y _06247_/X _06217_/A _06255_/X vssd1 vssd1 vccd1 vccd1 _13273_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_191_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06187_ _06032_/Y _06033_/Y _06035_/B _06186_/X vssd1 vssd1 vccd1 vccd1 _06187_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09946_ _08787_/Y _09943_/X _06255_/X _09938_/X _09941_/X vssd1 vssd1 vccd1 vccd1
+ _09946_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_104_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09877_ _09877_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09877_/X sky130_fd_sc_hd__or2_1
XFILLER_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08828_ _08836_/A vssd1 vssd1 vccd1 vccd1 _08828_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _12680_/Q vssd1 vssd1 vccd1 vccd1 _08759_/Y sky130_fd_sc_hd__inv_2
XPHY_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11769_/X _12111_/X _11774_/S vssd1 vssd1 vccd1 vccd1 _12432_/D sky130_fd_sc_hd__mux2_1
XPHY_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _13245_/Q _10738_/A _10779_/A _10717_/X _06430_/X vssd1 vssd1 vccd1 vccd1
+ _11139_/A sky130_fd_sc_hd__o221a_1
XPHY_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10652_ _11907_/X vssd1 vssd1 vccd1 vccd1 _10652_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10583_ _10583_/A _11386_/X vssd1 vssd1 vccd1 vccd1 _10583_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_186_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12322_ _12517_/CLK _12322_/D vssd1 vssd1 vccd1 vccd1 _12322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12253_ _12781_/Q _12854_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12253_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11204_ vssd1 vssd1 vccd1 vccd1 _11204_/HI _11204_/LO sky130_fd_sc_hd__conb_1
XFILLER_181_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12184_ _10702_/X _07020_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12184_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11135_ _11135_/A vssd1 vssd1 vccd1 vccd1 _11135_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11066_ _10773_/X _11037_/X _06386_/X _11058_/X _11038_/X vssd1 vssd1 vccd1 vccd1
+ _11066_/X sky130_fd_sc_hd__a221o_1
XFILLER_27_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10017_ _12622_/Q vssd1 vssd1 vccd1 vccd1 _10017_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11968_ _09297_/Y _09301_/Y _11969_/S vssd1 vssd1 vccd1 vccd1 _11968_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10919_ _12342_/Q vssd1 vssd1 vccd1 vccd1 _10919_/Y sky130_fd_sc_hd__inv_2
X_11899_ _10744_/Y _06583_/A _12760_/Q vssd1 vssd1 vccd1 vccd1 _11899_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06110_ _12722_/Q _12690_/Q _06109_/X vssd1 vssd1 vccd1 vccd1 _06175_/B sky130_fd_sc_hd__o21ai_1
XFILLER_117_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07090_ _11964_/S vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__inv_2
XFILLER_173_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06041_ _12741_/Q vssd1 vssd1 vccd1 vccd1 _06041_/Y sky130_fd_sc_hd__inv_2
Xoutput503 _11252_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput514 _11262_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__clkbuf_2
Xoutput525 _11272_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput536 _11282_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput547 _11292_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput558 _11302_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__clkbuf_2
Xoutput569 _11312_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09800_ _09800_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09800_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07992_ _08004_/A vssd1 vssd1 vccd1 vccd1 _07992_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09731_ _09747_/B vssd1 vssd1 vccd1 vccd1 _09731_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06943_ _13181_/Q vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__inv_2
XFILLER_28_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09662_ _13161_/Q _09475_/X _09649_/Y _09919_/B _09661_/X vssd1 vssd1 vccd1 vccd1
+ _09662_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_28_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06874_ _12039_/X _06872_/B _06872_/X vssd1 vssd1 vccd1 vccd1 _06874_/X sky130_fd_sc_hd__a21bo_1
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08613_ _08623_/A vssd1 vssd1 vccd1 vccd1 _08613_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09593_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09593_/X sky130_fd_sc_hd__or2_1
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08544_ _07069_/A _07074_/X _12752_/Q _12753_/Q _07042_/A vssd1 vssd1 vccd1 vccd1
+ _12753_/D sky130_fd_sc_hd__a32o_1
XPHY_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08475_ _13047_/Q vssd1 vssd1 vccd1 vccd1 _08475_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07426_ _07428_/A vssd1 vssd1 vccd1 vccd1 _07426_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07357_ _11436_/X _07353_/X _13060_/Q _07354_/X vssd1 vssd1 vccd1 vccd1 _13060_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06308_ _06313_/A vssd1 vssd1 vccd1 vccd1 _06308_/X sky130_fd_sc_hd__clkbuf_1
X_07288_ hold1/A _07285_/X _07287_/X _11514_/S vssd1 vssd1 vccd1 vccd1 _13081_/D sky130_fd_sc_hd__a22o_1
XFILLER_156_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09027_ _09288_/B _09027_/B vssd1 vssd1 vccd1 vccd1 _09027_/Y sky130_fd_sc_hd__nor2_1
X_06239_ _06245_/A vssd1 vssd1 vccd1 vccd1 _06239_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09929_ _12889_/Q _09935_/B vssd1 vssd1 vccd1 vccd1 _09929_/X sky130_fd_sc_hd__or2_1
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12940_ _12975_/CLK _12940_/D vssd1 vssd1 vccd1 vccd1 _12940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _12871_/CLK _12871_/D _08036_/X vssd1 vssd1 vccd1 vccd1 _12871_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _09899_/Y _12847_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__mux2_1
XPHY_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _11376_/X _11752_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11753_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10704_ _12761_/Q _12760_/Q vssd1 vssd1 vccd1 vccd1 _10704_/Y sky130_fd_sc_hd__nor2_2
XPHY_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _11683_/X _11377_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12384_/D sky130_fd_sc_hd__mux2_1
XPHY_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10635_ _11891_/X _10649_/B vssd1 vssd1 vccd1 vccd1 _10635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_186_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10566_ _12395_/D _12396_/D _10521_/A _09411_/Y _11390_/S vssd1 vssd1 vccd1 vccd1
+ _10566_/X sky130_fd_sc_hd__o221a_1
XFILLER_154_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12305_ _12939_/CLK _12965_/Q vssd1 vssd1 vccd1 vccd1 _12305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13285_ _13286_/CLK _13285_/D _06214_/A vssd1 vssd1 vccd1 vccd1 _13285_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10497_ _12502_/Q _09141_/B _09142_/B vssd1 vssd1 vccd1 vccd1 _10497_/X sky130_fd_sc_hd__a21bo_1
XFILLER_142_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12236_ _12235_/X _12638_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12236_/X sky130_fd_sc_hd__mux2_2
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12167_ _12168_/A0 _10488_/Y hold1/A vssd1 vssd1 vccd1 vccd1 _12167_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11118_ _10773_/A _11077_/X _13246_/Q _11086_/X _11087_/X vssd1 vssd1 vccd1 vccd1
+ _11118_/X sky130_fd_sc_hd__a221o_1
XFILLER_111_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12098_ _12429_/Q _10666_/Y _12141_/S vssd1 vssd1 vccd1 vccd1 _12098_/X sky130_fd_sc_hd__mux2_1
X_11049_ _11049_/A vssd1 vssd1 vccd1 vccd1 _11049_/Y sky130_fd_sc_hd__inv_2
Xinput7 io_in[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
XFILLER_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06590_ _12202_/X _12201_/X _12202_/X _12201_/X vssd1 vssd1 vccd1 vccd1 _06590_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08260_ _08282_/A vssd1 vssd1 vccd1 vccd1 _08260_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07211_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07211_/X sky130_fd_sc_hd__clkbuf_1
X_08191_ _08132_/X _08163_/X _08191_/C _08191_/D vssd1 vssd1 vccd1 vccd1 _08191_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_119_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07142_ _07152_/A vssd1 vssd1 vccd1 vccd1 _07142_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07073_ _07078_/A vssd1 vssd1 vccd1 vccd1 _07073_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06024_ _12749_/Q _12717_/Q vssd1 vssd1 vccd1 vccd1 _06025_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput377 _11163_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__clkbuf_2
Xoutput388 _11173_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput399 _11344_/X vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07975_ _07975_/A vssd1 vssd1 vccd1 vccd1 _07975_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ _09714_/A _09748_/A _09714_/C vssd1 vssd1 vccd1 vccd1 _09717_/A sky130_fd_sc_hd__or3_4
X_06926_ _11995_/X _06924_/B _06924_/X vssd1 vssd1 vccd1 vccd1 _06926_/X sky130_fd_sc_hd__a21bo_1
XFILLER_28_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ _09673_/A vssd1 vssd1 vccd1 vccd1 _09646_/B sky130_fd_sc_hd__inv_2
X_06857_ _06857_/A _06857_/B vssd1 vssd1 vccd1 vccd1 _06857_/Y sky130_fd_sc_hd__nor2_2
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09576_ _09576_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09576_/Y sky130_fd_sc_hd__nor2_2
XFILLER_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06788_ _12016_/X _12012_/X _12016_/X _12012_/X vssd1 vssd1 vccd1 vccd1 _06788_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_128_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08527_ _08519_/X _12242_/X _08514_/X _12758_/Q vssd1 vssd1 vccd1 vccd1 _12758_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_1_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08458_ _13064_/Q _10380_/B _12836_/Q vssd1 vssd1 vccd1 vccd1 _08474_/A sky130_fd_sc_hd__o21ai_1
XPHY_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07409_ _07409_/A _09976_/B _09295_/A vssd1 vssd1 vccd1 vccd1 _07409_/Y sky130_fd_sc_hd__nor3_4
XFILLER_184_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08389_ _08405_/A vssd1 vssd1 vccd1 vccd1 _08389_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10420_ _10420_/A _10420_/B vssd1 vssd1 vccd1 vccd1 _10422_/B sky130_fd_sc_hd__nor2_2
XFILLER_164_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10351_ _07839_/X _10352_/C _12905_/Q _10349_/B _10350_/X vssd1 vssd1 vccd1 vccd1
+ _10351_/X sky130_fd_sc_hd__o221a_1
XFILLER_152_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13070_ _12165_/X _13070_/D _07330_/X vssd1 vssd1 vccd1 vccd1 _13070_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10282_ _10280_/Y _10032_/X _10281_/Y _10028_/X vssd1 vssd1 vccd1 vccd1 _10282_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12021_ _11082_/X _11074_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _12021_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12923_ _12166_/X _12923_/D _07895_/X vssd1 vssd1 vccd1 vccd1 _12923_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12854_ _12868_/CLK _12854_/D _08081_/X vssd1 vssd1 vccd1 vccd1 _12854_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _09180_/B _11804_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11805_/X sky130_fd_sc_hd__mux2_1
XPHY_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _12888_/CLK _12785_/D _08408_/X vssd1 vssd1 vccd1 vccd1 _12785_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _09180_/C _11735_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11736_/X sky130_fd_sc_hd__mux2_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11667_ _11379_/X _09186_/B _11675_/S vssd1 vssd1 vccd1 vccd1 _11667_/X sky130_fd_sc_hd__mux2_1
XPHY_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10618_ _12411_/D _12412_/D _10619_/B _10617_/Y vssd1 vssd1 vccd1 vccd1 _10618_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11598_ _10458_/Y _09180_/C _11603_/S vssd1 vssd1 vccd1 vccd1 _11598_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10549_ _09331_/A _09331_/B _10548_/Y vssd1 vssd1 vccd1 vccd1 _10549_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13268_ _13268_/CLK _13268_/D _06280_/X vssd1 vssd1 vccd1 vccd1 _13268_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12219_ _06311_/Y _13155_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__mux2_1
X_13199_ _13201_/CLK _13199_/D _06780_/X vssd1 vssd1 vccd1 vccd1 _13199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07760_ _12586_/Q _07760_/B vssd1 vssd1 vccd1 vccd1 _07761_/B sky130_fd_sc_hd__or2_1
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06711_ _06699_/X _06703_/X _06704_/X vssd1 vssd1 vccd1 vccd1 _06711_/X sky130_fd_sc_hd__a21bo_1
XFILLER_65_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07691_ _07686_/B _07690_/Y _07672_/C _12307_/Q vssd1 vssd1 vccd1 vccd1 _07717_/A
+ sky130_fd_sc_hd__o31a_2
X_09430_ _09379_/Y _12408_/D _12546_/Q _09428_/Y _09429_/X vssd1 vssd1 vccd1 vccd1
+ _09430_/X sky130_fd_sc_hd__o221a_1
X_06642_ _11901_/X _12196_/X _11901_/X _12196_/X vssd1 vssd1 vccd1 vccd1 _06642_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_25_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _09341_/Y _12410_/Q _12466_/Q _09342_/Y _09360_/X vssd1 vssd1 vccd1 vccd1
+ _09371_/B sky130_fd_sc_hd__o221a_1
XFILLER_178_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06573_ _06573_/A _06573_/B vssd1 vssd1 vccd1 vccd1 _06573_/Y sky130_fd_sc_hd__nor2_2
XFILLER_127_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12490_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08312_ _12822_/Q _11597_/X _08321_/S vssd1 vssd1 vccd1 vccd1 _12822_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09292_ _09269_/X _09292_/B vssd1 vssd1 vccd1 vccd1 _12302_/D sky130_fd_sc_hd__nand2b_1
XFILLER_127_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08243_ _13098_/Q _10449_/B _13101_/Q _10454_/A _08242_/X vssd1 vssd1 vccd1 vccd1
+ _08246_/C sky130_fd_sc_hd__o221a_1
XFILLER_166_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08174_ _08116_/Y _08117_/X _13145_/Q _08122_/Y _08173_/Y vssd1 vssd1 vccd1 vccd1
+ _08175_/D sky130_fd_sc_hd__o221a_1
XFILLER_180_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07125_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07125_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07056_ _07053_/X _07040_/X _06300_/Y _13157_/Q _07042_/X vssd1 vssd1 vccd1 vccd1
+ _13157_/D sky130_fd_sc_hd__a32o_1
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06007_ _11969_/S _11964_/S vssd1 vssd1 vccd1 vccd1 _09981_/C sky130_fd_sc_hd__or2_2
XFILLER_121_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07958_ _12897_/Q _11486_/X _07962_/S vssd1 vssd1 vccd1 vccd1 _12897_/D sky130_fd_sc_hd__mux2_1
X_06909_ _13185_/Q vssd1 vssd1 vccd1 vccd1 _06909_/Y sky130_fd_sc_hd__inv_2
X_07889_ _12836_/Q vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__inv_2
XFILLER_29_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09628_ _09471_/X _09624_/X _09625_/Y _09627_/X vssd1 vssd1 vccd1 vccd1 _09628_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_83_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09559_ _09952_/A _09949_/A _09572_/A _09558_/B _09566_/B vssd1 vssd1 vccd1 vccd1
+ _09559_/X sky130_fd_sc_hd__a221o_1
XFILLER_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12570_ _12570_/CLK _12570_/D vssd1 vssd1 vccd1 vccd1 _12570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ _12810_/Q input357/X _11522_/S vssd1 vssd1 vccd1 vccd1 _11521_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11452_ _12895_/Q _09185_/C _11459_/S vssd1 vssd1 vccd1 vccd1 _11452_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10403_ _10411_/A vssd1 vssd1 vccd1 vccd1 _10458_/A sky130_fd_sc_hd__clkbuf_4
X_11383_ _10566_/X _12396_/D _11392_/S vssd1 vssd1 vccd1 vccd1 _11383_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10334_ _10333_/A _10333_/B _10335_/B _10324_/A vssd1 vssd1 vccd1 vccd1 _10334_/Y
+ sky130_fd_sc_hd__a211oi_4
X_13122_ _12168_/X _13122_/D _07173_/X vssd1 vssd1 vccd1 vccd1 _13122_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13053_ _12165_/X _13053_/D _07373_/X vssd1 vssd1 vccd1 vccd1 _13053_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10265_ _10263_/Y _10032_/X _10264_/Y _10028_/X vssd1 vssd1 vccd1 vccd1 _10265_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12004_ _11106_/X _11098_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12004_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10196_ _12853_/Q vssd1 vssd1 vccd1 vccd1 _10196_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12906_ _12166_/X _12906_/D _07934_/X vssd1 vssd1 vccd1 vccd1 _12906_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12837_ _12166_/A0 _12837_/D _08264_/X vssd1 vssd1 vccd1 vccd1 _12837_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12769_/CLK _12768_/D _08501_/X vssd1 vssd1 vccd1 vccd1 _12768_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11719_ _10652_/Y _10653_/Y _11818_/S vssd1 vssd1 vccd1 vccd1 _11719_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12699_ _12717_/CLK _12699_/D _08706_/X vssd1 vssd1 vccd1 vccd1 _12699_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput10 io_in[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
Xinput21 io_in[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_1
Xinput32 io_in[3] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_2
Xinput43 la_data_in[103] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_1
XFILLER_174_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput54 la_data_in[113] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_1
XFILLER_190_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput65 la_data_in[123] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_1
Xinput76 la_data_in[18] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__buf_1
XFILLER_116_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput87 la_data_in[28] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__buf_1
Xinput98 la_data_in[38] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__buf_1
XFILLER_66_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_137_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12753_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_104_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ _08930_/A _10643_/A vssd1 vssd1 vccd1 vccd1 _08931_/A sky130_fd_sc_hd__or2_2
XFILLER_112_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08861_ _08849_/X _06323_/Y _08852_/X _12644_/Q vssd1 vssd1 vccd1 vccd1 _12644_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_112_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater611 _11831_/S vssd1 vssd1 vccd1 vccd1 _11851_/S sky130_fd_sc_hd__buf_8
X_07812_ _13015_/Q _10333_/A _07808_/Y _12903_/Q _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07819_/C sky130_fd_sc_hd__a221o_1
XFILLER_96_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08792_ _08839_/A vssd1 vssd1 vccd1 vccd1 _08807_/A sky130_fd_sc_hd__clkbuf_2
Xrepeater622 _11433_/S vssd1 vssd1 vccd1 vccd1 _11443_/S sky130_fd_sc_hd__buf_4
XFILLER_42_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater633 input358/X vssd1 vssd1 vccd1 vccd1 _09185_/A sky130_fd_sc_hd__buf_8
Xrepeater644 input337/X vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__buf_8
X_07743_ _12943_/Q _07740_/Y _07750_/B _09282_/B vssd1 vssd1 vccd1 vccd1 _12943_/D
+ sky130_fd_sc_hd__o22a_1
X_07674_ _09276_/C vssd1 vssd1 vccd1 vccd1 _09279_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09413_ _12454_/Q _10586_/A _12542_/Q _10611_/A vssd1 vssd1 vccd1 vccd1 _09413_/X
+ sky130_fd_sc_hd__a22o_1
X_06625_ _06625_/A _06625_/B vssd1 vssd1 vccd1 vccd1 _06625_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09344_ _09343_/Y _12403_/Q _09343_/Y _12403_/Q vssd1 vssd1 vccd1 vccd1 _09344_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_34_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06556_ _12621_/Q vssd1 vssd1 vccd1 vccd1 _06556_/X sky130_fd_sc_hd__buf_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09275_ _09269_/A _12303_/Q _09271_/C _09271_/X _09274_/Y vssd1 vssd1 vccd1 vccd1
+ _09277_/C sky130_fd_sc_hd__a311o_1
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06487_ _06522_/A vssd1 vssd1 vccd1 vccd1 _06487_/X sky130_fd_sc_hd__clkbuf_1
X_08226_ _13083_/Q vssd1 vssd1 vccd1 vccd1 _08226_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08157_ _12815_/Q vssd1 vssd1 vccd1 vccd1 _10433_/A sky130_fd_sc_hd__inv_2
XFILLER_180_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07108_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07108_/X sky130_fd_sc_hd__clkbuf_1
X_08088_ _08098_/A vssd1 vssd1 vccd1 vccd1 _08088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07039_ _07059_/A vssd1 vssd1 vccd1 vccd1 _07074_/A sky130_fd_sc_hd__inv_2
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10050_ _10113_/A vssd1 vssd1 vccd1 vccd1 _10277_/A sky130_fd_sc_hd__inv_2
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10952_ _12534_/Q vssd1 vssd1 vccd1 vccd1 _10952_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10883_ _10888_/C _10882_/Y _10888_/C _10882_/Y vssd1 vssd1 vccd1 vccd1 _12336_/D
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_32_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12622_ _13154_/CLK _12622_/D _08915_/X vssd1 vssd1 vccd1 vccd1 _12622_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ _13154_/CLK _12553_/D _09065_/X vssd1 vssd1 vccd1 vccd1 _12553_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11504_ _10379_/X _09179_/D _11513_/S vssd1 vssd1 vccd1 vccd1 _11504_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12484_ _12168_/A0 _12484_/D vssd1 vssd1 vccd1 vccd1 _12484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ _12910_/Q _09179_/A _11443_/S vssd1 vssd1 vccd1 vccd1 _11435_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11366_ _11365_/X _12444_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11366_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10317_ _12893_/Q _10371_/A vssd1 vssd1 vccd1 vccd1 _10317_/Y sky130_fd_sc_hd__nor2_1
X_13105_ _12167_/X _13105_/D _07224_/X vssd1 vssd1 vccd1 vccd1 _13105_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11297_ vssd1 vssd1 vccd1 vccd1 _11297_/HI _11297_/LO sky130_fd_sc_hd__conb_1
XFILLER_152_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10248_ _13266_/Q vssd1 vssd1 vccd1 vccd1 _10248_/Y sky130_fd_sc_hd__inv_2
X_13036_ _12164_/X _13036_/D _07424_/X vssd1 vssd1 vccd1 vccd1 _13036_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10179_ _12852_/Q vssd1 vssd1 vccd1 vccd1 _10179_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06410_ _13239_/Q vssd1 vssd1 vccd1 vccd1 _06410_/X sky130_fd_sc_hd__buf_2
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07390_ _11423_/X _07384_/X _13047_/Q _07385_/X vssd1 vssd1 vccd1 vccd1 _13047_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06341_ _06339_/X _06340_/X _06339_/X _06340_/X vssd1 vssd1 vccd1 vccd1 _06342_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_188_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ _10227_/A _12147_/X vssd1 vssd1 vccd1 vccd1 _12558_/D sky130_fd_sc_hd__nor2b_4
XFILLER_8_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06272_ _06272_/A vssd1 vssd1 vccd1 vccd1 _06306_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_191_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08011_ _12881_/Q _07996_/X _07296_/X _07998_/X vssd1 vssd1 vccd1 vccd1 _12881_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09962_ _08739_/Y _09897_/A _11963_/S _09892_/A _09941_/A vssd1 vssd1 vccd1 vccd1
+ _09962_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_98_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08913_ _08898_/A _06346_/Y _08908_/X _12623_/Q vssd1 vssd1 vccd1 vccd1 _12623_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_83_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09893_ _09939_/B vssd1 vssd1 vccd1 vccd1 _09910_/B sky130_fd_sc_hd__buf_1
XFILLER_58_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08844_ _08851_/A vssd1 vssd1 vccd1 vccd1 _08844_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08775_ _08774_/Y _08760_/X _06233_/X _08764_/X vssd1 vssd1 vccd1 vccd1 _12676_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12410_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07726_ _07726_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07726_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07657_ _07678_/A _12946_/Q _12948_/Q _07657_/D vssd1 vssd1 vccd1 vccd1 _07658_/C
+ sky130_fd_sc_hd__or4_4
XPHY_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06608_ _06769_/A vssd1 vssd1 vccd1 vccd1 _06608_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_186_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07588_ _09269_/A vssd1 vssd1 vccd1 vccd1 _09284_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09327_ _09327_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09328_/B sky130_fd_sc_hd__or2_1
XFILLER_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06539_ _12172_/X _11135_/A vssd1 vssd1 vccd1 vccd1 _06539_/X sky130_fd_sc_hd__or2_1
XFILLER_159_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09258_ _12451_/Q _09251_/A _09242_/A _09083_/A vssd1 vssd1 vccd1 vccd1 _12451_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08209_ _08209_/A _08209_/B _08209_/C _08208_/X vssd1 vssd1 vccd1 vccd1 _08247_/A
+ sky130_fd_sc_hd__or4b_4
X_09189_ _10655_/B _11817_/S vssd1 vssd1 vccd1 vccd1 _09215_/A sky130_fd_sc_hd__or2_4
XFILLER_147_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11220_ vssd1 vssd1 vccd1 vccd1 _11220_/HI _11220_/LO sky130_fd_sc_hd__conb_1
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11151_ vssd1 vssd1 vccd1 vccd1 _11151_/HI _11151_/LO sky130_fd_sc_hd__conb_1
XFILLER_150_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10102_ _10101_/Y _10137_/A _09900_/Y _10003_/A vssd1 vssd1 vccd1 vccd1 _10107_/C
+ sky130_fd_sc_hd__o22a_1
X_11082_ _10773_/X _11054_/X _06386_/X _11055_/X _11060_/X vssd1 vssd1 vccd1 vccd1
+ _11082_/X sky130_fd_sc_hd__a221o_1
Xinput200 la_oenb[14] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__buf_1
Xinput211 la_oenb[24] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__buf_1
Xinput222 la_oenb[34] vssd1 vssd1 vccd1 vccd1 input222/X sky130_fd_sc_hd__buf_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10033_ _10141_/A vssd1 vssd1 vccd1 vccd1 _10033_/X sky130_fd_sc_hd__clkbuf_2
Xinput233 la_oenb[44] vssd1 vssd1 vccd1 vccd1 input233/X sky130_fd_sc_hd__buf_1
XFILLER_49_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput244 la_oenb[54] vssd1 vssd1 vccd1 vccd1 input244/X sky130_fd_sc_hd__buf_1
Xinput255 la_oenb[64] vssd1 vssd1 vccd1 vccd1 input255/X sky130_fd_sc_hd__buf_1
XFILLER_102_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput266 la_oenb[74] vssd1 vssd1 vccd1 vccd1 input266/X sky130_fd_sc_hd__buf_1
XFILLER_102_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput277 la_oenb[84] vssd1 vssd1 vccd1 vccd1 input277/X sky130_fd_sc_hd__buf_1
Xinput288 la_oenb[94] vssd1 vssd1 vccd1 vccd1 input288/X sky130_fd_sc_hd__buf_1
XFILLER_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput299 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 _09071_/D sky130_fd_sc_hd__buf_1
XFILLER_63_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11984_ _09434_/C _09434_/X _12549_/Q vssd1 vssd1 vccd1 vccd1 _12550_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10935_ _10934_/A _10933_/Y _10947_/B _10933_/A vssd1 vssd1 vccd1 vccd1 _12343_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10866_ _12518_/Q _12330_/Q _10843_/Y vssd1 vssd1 vccd1 vccd1 _10866_/X sky130_fd_sc_hd__a21o_1
X_12605_ _13008_/CLK _12605_/D vssd1 vssd1 vccd1 vccd1 _12605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10797_ _12510_/Q vssd1 vssd1 vccd1 vccd1 _10799_/A sky130_fd_sc_hd__inv_2
XFILLER_185_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12536_ _12541_/CLK _12536_/D vssd1 vssd1 vccd1 vccd1 _12536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12467_ _12467_/CLK _12467_/D vssd1 vssd1 vccd1 vccd1 _12467_/Q sky130_fd_sc_hd__dfxtp_1
X_11418_ _12893_/Q _09184_/A _11449_/S vssd1 vssd1 vccd1 vccd1 _11418_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12398_ _12415_/CLK _12398_/D vssd1 vssd1 vccd1 vccd1 _12398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11349_ _09446_/X _12986_/Q _11356_/S vssd1 vssd1 vccd1 vccd1 _12313_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13019_ _12164_/X _13019_/D _07467_/X vssd1 vssd1 vccd1 vccd1 _13019_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_67_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06890_ _06890_/A _06890_/B vssd1 vssd1 vccd1 vccd1 _06890_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08560_ _08569_/A vssd1 vssd1 vccd1 vccd1 _08560_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07511_ _09186_/A vssd1 vssd1 vccd1 vccd1 _09227_/A sky130_fd_sc_hd__inv_2
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08491_ _13054_/Q _07839_/X _13054_/Q _07839_/X vssd1 vssd1 vccd1 vccd1 _08491_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07442_ _11470_/X _07429_/X _13029_/Q _07430_/X vssd1 vssd1 vccd1 vccd1 _13029_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07373_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07373_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09112_ _12526_/Q _09107_/X input336/X _09108_/X vssd1 vssd1 vccd1 vccd1 _12526_/D
+ sky130_fd_sc_hd__a22o_1
X_06324_ _06303_/X _06314_/X _06323_/Y _13261_/Q _06306_/X vssd1 vssd1 vccd1 vccd1
+ _13261_/D sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_152_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13257_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09043_ _09043_/A _09043_/B _09043_/C _09433_/B vssd1 vssd1 vccd1 vccd1 _10190_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_159_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06255_ _06060_/A _06254_/X _06060_/A _06254_/X vssd1 vssd1 vccd1 vccd1 _06255_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_163_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06186_ _06185_/A _06171_/X _06184_/X _06185_/X _06154_/A vssd1 vssd1 vccd1 vccd1
+ _06186_/X sky130_fd_sc_hd__o221a_1
XFILLER_117_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09945_ _08790_/Y _09943_/X _06260_/X _09938_/X _09941_/X vssd1 vssd1 vccd1 vccd1
+ _09945_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_131_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09876_ _09877_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09876_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08827_ _08814_/X _08817_/X _06332_/Y _12658_/Q _08567_/A vssd1 vssd1 vccd1 vccd1
+ _12658_/D sky130_fd_sc_hd__a32o_1
XFILLER_45_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _08769_/A vssd1 vssd1 vccd1 vccd1 _08758_/X sky130_fd_sc_hd__clkbuf_1
XPHY_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _12956_/Q _07707_/X _12955_/Q _07705_/X _07703_/X vssd1 vssd1 vccd1 vccd1
+ _12956_/D sky130_fd_sc_hd__o221a_1
XPHY_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _08699_/A vssd1 vssd1 vccd1 vccd1 _08689_/X sky130_fd_sc_hd__clkbuf_1
XPHY_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ _13245_/Q vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__inv_2
XFILLER_81_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10651_ _12424_/Q _08932_/B _10650_/Y _08931_/A vssd1 vssd1 vccd1 vccd1 _10651_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10582_ _12401_/D _09415_/Y _10578_/Y _12402_/D _10579_/X vssd1 vssd1 vccd1 vccd1
+ _10582_/X sky130_fd_sc_hd__a32o_1
XFILLER_155_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12321_ _12577_/CLK _12321_/D vssd1 vssd1 vccd1 vccd1 _12321_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_154_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12252_ _12251_/X _12646_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12252_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11203_ vssd1 vssd1 vccd1 vccd1 _11203_/HI _11203_/LO sky130_fd_sc_hd__conb_1
XFILLER_108_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12183_ _10697_/X _10694_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _12183_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11134_ _10767_/A _10788_/X _13247_/Q _11111_/X _11112_/X vssd1 vssd1 vccd1 vccd1
+ _11134_/X sky130_fd_sc_hd__a221o_1
XFILLER_150_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11065_ _06379_/X _11045_/X _11032_/X _10763_/X _11034_/X vssd1 vssd1 vccd1 vccd1
+ _11065_/X sky130_fd_sc_hd__a32o_1
XFILLER_62_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10016_ _09284_/B _10015_/Y _12303_/Q _11971_/X vssd1 vssd1 vccd1 vccd1 _10016_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11967_ _09300_/Y _09302_/Y _11967_/S vssd1 vssd1 vccd1 vccd1 _11967_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10918_ _12530_/Q vssd1 vssd1 vccd1 vccd1 _10918_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11898_ _06586_/A _10748_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__mux2_2
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10849_ _12520_/Q vssd1 vssd1 vccd1 vccd1 _10849_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12519_ _12801_/CLK _12519_/D vssd1 vssd1 vccd1 vccd1 _12519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_172_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06040_ _12743_/Q _12711_/Q _06038_/Y _06039_/Y vssd1 vssd1 vccd1 vccd1 _06046_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput504 _11253_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__clkbuf_2
XFILLER_172_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput515 _11263_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput526 _11273_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
Xoutput537 _11283_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__clkbuf_2
Xoutput548 _11293_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__clkbuf_2
Xoutput559 _11303_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07991_ _12888_/Q _07974_/X _07990_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _12888_/D
+ sky130_fd_sc_hd__a22o_1
X_09730_ _09709_/A _09729_/A _09709_/Y _09729_/Y vssd1 vssd1 vccd1 vccd1 _09747_/B
+ sky130_fd_sc_hd__o22a_1
X_06942_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06942_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09661_ _09673_/B _09659_/X _09660_/Y vssd1 vssd1 vccd1 vccd1 _09661_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06873_ _11997_/X _11994_/X _06872_/X vssd1 vssd1 vccd1 vccd1 _06873_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08612_ _08642_/A vssd1 vssd1 vccd1 vccd1 _08623_/A sky130_fd_sc_hd__clkbuf_2
X_09592_ _09592_/A _09592_/B vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__or2_1
XFILLER_94_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08543_ _08569_/A vssd1 vssd1 vccd1 vccd1 _08543_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08474_ _08474_/A _08474_/B _08474_/C _08473_/X vssd1 vssd1 vccd1 vccd1 _08474_/X
+ sky130_fd_sc_hd__or4b_4
XPHY_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07425_ _11477_/X _07412_/X _13036_/Q _07415_/X vssd1 vssd1 vccd1 vccd1 _13036_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07356_ _07360_/A vssd1 vssd1 vccd1 vccd1 _07356_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06307_ _06303_/X _06281_/X _06305_/X _13264_/Q _06306_/X vssd1 vssd1 vccd1 vccd1
+ _13264_/D sky130_fd_sc_hd__a32o_1
XFILLER_109_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07287_ _09242_/A vssd1 vssd1 vccd1 vccd1 _07287_/X sky130_fd_sc_hd__buf_2
XFILLER_109_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ _10015_/B _12302_/Q vssd1 vssd1 vccd1 vccd1 _09027_/B sky130_fd_sc_hd__nand2_2
X_06238_ _06236_/Y _06216_/X _06217_/X _06237_/X vssd1 vssd1 vccd1 vccd1 _13276_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_145_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06169_ _13285_/Q vssd1 vssd1 vccd1 vccd1 _06169_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09928_ _12666_/Q vssd1 vssd1 vccd1 vccd1 _09928_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09859_ _09860_/A _09866_/B vssd1 vssd1 vccd1 vccd1 _09859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12870_ _12870_/CLK _12870_/D _08039_/X vssd1 vssd1 vccd1 vccd1 _12870_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11821_ _09895_/Y _12846_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11821_/X sky130_fd_sc_hd__mux2_1
XPHY_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _09186_/B _11751_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11752_/X sky130_fd_sc_hd__mux2_1
XPHY_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _13240_/Q _07019_/A _10693_/X _11071_/A _06637_/Y vssd1 vssd1 vccd1 vccd1
+ _11036_/A sky130_fd_sc_hd__o221a_1
XFILLER_186_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11377_/X _09244_/B _11691_/S vssd1 vssd1 vccd1 vccd1 _11683_/X sky130_fd_sc_hd__mux2_1
XPHY_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10634_ _11891_/X vssd1 vssd1 vccd1 vccd1 _10634_/Y sky130_fd_sc_hd__inv_2
XPHY_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10565_ _12395_/D _10570_/A vssd1 vssd1 vccd1 vccd1 _10565_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12304_ _12576_/CLK _12304_/D vssd1 vssd1 vccd1 vccd1 _12304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13284_ _13286_/CLK _13284_/D _06190_/X vssd1 vssd1 vccd1 vccd1 _13284_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10496_ _12501_/Q _09140_/B _09141_/B vssd1 vssd1 vccd1 vccd1 _10496_/X sky130_fd_sc_hd__a21bo_1
XFILLER_120_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12235_ _12772_/Q _12845_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12235_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12166_ _12166_/A0 _07887_/X _12837_/Q vssd1 vssd1 vccd1 vccd1 _12166_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11117_ _10763_/X _11075_/X _13248_/Q _11083_/X _11084_/X vssd1 vssd1 vccd1 vccd1
+ _11117_/X sky130_fd_sc_hd__a221o_1
XFILLER_7_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12097_ _06446_/B _10710_/Y _12768_/Q vssd1 vssd1 vccd1 vccd1 _12199_/S sky130_fd_sc_hd__mux2_8
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11048_ _10696_/X _10746_/X _06404_/X _07008_/X _10747_/X vssd1 vssd1 vccd1 vccd1
+ _11048_/X sky130_fd_sc_hd__a221o_1
Xinput8 io_in[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_1
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12999_ _12999_/CLK _12999_/D vssd1 vssd1 vccd1 vccd1 _12999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07210_ _11576_/X _07201_/X _13111_/Q _07204_/X vssd1 vssd1 vccd1 vccd1 _13111_/D
+ sky130_fd_sc_hd__a22o_1
X_08190_ _08179_/X _08190_/B _08190_/C _08190_/D vssd1 vssd1 vccd1 vccd1 _08191_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_119_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07141_ _11536_/X _07130_/X _13135_/Q _07131_/X vssd1 vssd1 vccd1 vccd1 _13135_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07072_ _07069_/X _07058_/X _06332_/Y _13151_/Q _07059_/X vssd1 vssd1 vccd1 vccd1
+ _13151_/D sky130_fd_sc_hd__a32o_1
XFILLER_69_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06023_ _12749_/Q _12717_/Q vssd1 vssd1 vccd1 vccd1 _06025_/A sky130_fd_sc_hd__and2_1
XFILLER_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput367 _11148_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput378 _11149_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__clkbuf_2
Xoutput389 _11154_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07974_ _07996_/A vssd1 vssd1 vccd1 vccd1 _07974_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09713_ _09713_/A _09713_/B vssd1 vssd1 vccd1 vccd1 _09748_/A sky130_fd_sc_hd__or2_2
X_06925_ _12001_/X _11998_/X _06924_/X vssd1 vssd1 vccd1 vccd1 _06925_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09644_ _09643_/A _09643_/B _09659_/A vssd1 vssd1 vccd1 vccd1 _09673_/A sky130_fd_sc_hd__a21oi_2
X_06856_ _06864_/A _06864_/B vssd1 vssd1 vccd1 vccd1 _06857_/B sky130_fd_sc_hd__and2_1
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09575_ _09556_/Y _09574_/B _09609_/A _09574_/X vssd1 vssd1 vccd1 vccd1 _09582_/A
+ sky130_fd_sc_hd__o211ai_2
X_06787_ _12037_/X _06785_/B _06785_/X vssd1 vssd1 vccd1 vccd1 _06787_/X sky130_fd_sc_hd__a21bo_1
XFILLER_36_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08526_ _08533_/A vssd1 vssd1 vccd1 vccd1 _08526_/X sky130_fd_sc_hd__clkbuf_1
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08457_ _08457_/A _08457_/B _08457_/C _08456_/X vssd1 vssd1 vccd1 vccd1 _08457_/X
+ sky130_fd_sc_hd__or4b_4
XPHY_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07408_ _07408_/A vssd1 vssd1 vccd1 vccd1 _07408_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08388_ _08521_/A vssd1 vssd1 vccd1 vccd1 _08405_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07339_ _07369_/A vssd1 vssd1 vccd1 vccd1 _07339_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _10372_/A vssd1 vssd1 vccd1 vccd1 _10350_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09009_ _09009_/A vssd1 vssd1 vccd1 vccd1 _09016_/A sky130_fd_sc_hd__buf_1
X_10281_ _12858_/Q vssd1 vssd1 vccd1 vccd1 _10281_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12020_ _11067_/X _11061_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _12020_/X sky130_fd_sc_hd__mux2_2
XFILLER_105_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12922_ _12166_/X _12922_/D _07897_/X vssd1 vssd1 vccd1 vccd1 _12922_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12853_ _12868_/CLK _12853_/D _08085_/X vssd1 vssd1 vccd1 vccd1 _12853_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _12071_/X _12489_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11804_/X sky130_fd_sc_hd__mux2_1
XPHY_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12784_ _12942_/CLK _12784_/D _08410_/X vssd1 vssd1 vccd1 vccd1 _12784_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_199_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11367_/X _12488_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11735_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _11665_/X _11381_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12375_/D sky130_fd_sc_hd__mux2_1
XPHY_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10617_ _10617_/A vssd1 vssd1 vccd1 vccd1 _10617_/Y sky130_fd_sc_hd__inv_2
XPHY_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11597_ _10453_/X _09180_/D _11603_/S vssd1 vssd1 vccd1 vccd1 _11597_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10548_ _10548_/A vssd1 vssd1 vccd1 vccd1 _10548_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13267_ _13269_/CLK _13267_/D _06288_/X vssd1 vssd1 vccd1 vccd1 _13267_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10479_ _10477_/A _10477_/B _10474_/A _10478_/Y vssd1 vssd1 vccd1 vccd1 _10479_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_170_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12218_ _12217_/X _12629_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12218_/X sky130_fd_sc_hd__mux2_1
X_13198_ _13201_/CLK _13198_/D _06795_/X vssd1 vssd1 vccd1 vccd1 _13198_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12149_ _09998_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12149_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06710_ _13207_/Q vssd1 vssd1 vccd1 vccd1 _06710_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07690_ _07690_/A _07690_/B vssd1 vssd1 vccd1 vccd1 _07690_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06641_ _12198_/X _10765_/A _06639_/X vssd1 vssd1 vccd1 vccd1 _06641_/X sky130_fd_sc_hd__a21bo_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09360_ _12543_/Q _12412_/Q _12543_/Q _12412_/Q vssd1 vssd1 vccd1 vccd1 _09360_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_06572_ _06576_/A _06576_/B vssd1 vssd1 vccd1 vccd1 _06573_/B sky130_fd_sc_hd__and2_1
XFILLER_33_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08311_ _08311_/A vssd1 vssd1 vccd1 vccd1 _08311_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09291_ _13006_/Q _07512_/Y _09261_/X _09279_/B _09290_/X vssd1 vssd1 vccd1 vccd1
+ _09292_/B sky130_fd_sc_hd__o32a_1
XFILLER_61_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08242_ _13111_/Q _10482_/A _13095_/Q _10439_/A vssd1 vssd1 vccd1 vccd1 _08242_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_165_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_59_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12993_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_159_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08173_ _13130_/Q _10449_/B vssd1 vssd1 vccd1 vccd1 _08173_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07124_ _07154_/A vssd1 vssd1 vccd1 vccd1 _07137_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07055_ _07063_/A vssd1 vssd1 vccd1 vccd1 _07055_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06006_ _11966_/S vssd1 vssd1 vccd1 vccd1 _09986_/D sky130_fd_sc_hd__inv_2
XFILLER_114_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07957_ _07961_/A vssd1 vssd1 vccd1 vccd1 _07957_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06908_ _06916_/A vssd1 vssd1 vccd1 vccd1 _06908_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07888_ _07888_/A vssd1 vssd1 vccd1 vccd1 _07888_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ _09626_/Y _07735_/A _12873_/Q _12614_/Q vssd1 vssd1 vccd1 vccd1 _09627_/X
+ sky130_fd_sc_hd__a22o_1
X_06839_ _06863_/A vssd1 vssd1 vccd1 vccd1 _06839_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09558_ _09572_/A _09558_/B vssd1 vssd1 vccd1 vccd1 _09566_/B sky130_fd_sc_hd__nor2_1
XFILLER_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08509_ _08518_/A vssd1 vssd1 vccd1 vccd1 _08509_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_196_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09489_ _13168_/Q _09488_/X _13168_/Q _09488_/X vssd1 vssd1 vccd1 vccd1 _09490_/B
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ _12809_/Q _09185_/B _11522_/S vssd1 vssd1 vccd1 vccd1 _11520_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11451_ _12894_/Q _09185_/D _11459_/S vssd1 vssd1 vccd1 vccd1 _11451_/X sky130_fd_sc_hd__mux2_1
XPHY_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10402_ _13146_/Q _12554_/Q vssd1 vssd1 vccd1 vccd1 _10402_/X sky130_fd_sc_hd__or2_1
X_11382_ _10589_/Y _12403_/D _11404_/S vssd1 vssd1 vccd1 vccd1 _11382_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13121_ _12168_/X _13121_/D _07175_/X vssd1 vssd1 vccd1 vccd1 _13121_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10333_ _10333_/A _10333_/B vssd1 vssd1 vccd1 vccd1 _10335_/B sky130_fd_sc_hd__nor2_4
XFILLER_194_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13052_ _12165_/X _13052_/D _07375_/X vssd1 vssd1 vccd1 vccd1 _13052_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10264_ _12857_/Q vssd1 vssd1 vccd1 vccd1 _10264_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12003_ _11079_/Y _10768_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _12003_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10195_ _13263_/Q vssd1 vssd1 vccd1 vccd1 _10195_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12905_ _12166_/X _12905_/D _07937_/X vssd1 vssd1 vccd1 vccd1 _12905_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12836_ _12166_/A0 _12836_/D _08266_/X vssd1 vssd1 vccd1 vccd1 _12836_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12767_ _12769_/CLK _12767_/D _08503_/X vssd1 vssd1 vccd1 vccd1 _12767_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11718_ _11717_/X _10648_/Y _11774_/S vssd1 vssd1 vccd1 vccd1 _12423_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12698_ _12717_/CLK _12698_/D _08708_/X vssd1 vssd1 vccd1 vccd1 _12698_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_175_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput11 io_in[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_1
X_11649_ _10526_/Y _10529_/Y _11691_/S vssd1 vssd1 vccd1 vccd1 _11649_/X sky130_fd_sc_hd__mux2_1
Xinput22 io_in[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_1
XFILLER_156_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput33 io_in[4] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_1
XFILLER_190_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput44 la_data_in[104] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_1
Xinput55 la_data_in[114] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_1
Xinput66 la_data_in[124] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_1
XFILLER_122_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput77 la_data_in[19] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__buf_1
Xinput88 la_data_in[29] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__buf_1
XFILLER_116_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput99 la_data_in[39] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__buf_1
XFILLER_66_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08860_ _08866_/A vssd1 vssd1 vccd1 vccd1 _08860_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_123_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07811_ _13040_/Q _07809_/Y _13022_/Q _10352_/A vssd1 vssd1 vccd1 vccd1 _07811_/X
+ sky130_fd_sc_hd__a22o_1
Xrepeater612 _12103_/S vssd1 vssd1 vccd1 vccd1 _12142_/S sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_106_wb_clk_i _12726_/CLK vssd1 vssd1 vccd1 vccd1 _12725_/CLK sky130_fd_sc_hd__clkbuf_16
X_08791_ _08790_/Y _08781_/X _06260_/X _08764_/A vssd1 vssd1 vccd1 vccd1 _12671_/D
+ sky130_fd_sc_hd__o22ai_1
Xrepeater623 _11422_/S vssd1 vssd1 vccd1 vccd1 _11433_/S sky130_fd_sc_hd__buf_6
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater634 input357/X vssd1 vssd1 vccd1 vccd1 _09184_/B sky130_fd_sc_hd__buf_8
Xrepeater645 input336/X vssd1 vssd1 vccd1 vccd1 _09179_/B sky130_fd_sc_hd__buf_8
X_07742_ _08837_/A _07742_/B vssd1 vssd1 vccd1 vccd1 _09282_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07673_ _12307_/Q _07679_/A vssd1 vssd1 vccd1 vccd1 _07676_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09412_ _12411_/D vssd1 vssd1 vccd1 vccd1 _10611_/A sky130_fd_sc_hd__inv_2
X_06624_ _06650_/A vssd1 vssd1 vccd1 vccd1 _06624_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09343_ _12451_/Q vssd1 vssd1 vccd1 vccd1 _09343_/Y sky130_fd_sc_hd__inv_2
X_06555_ _06549_/Y _06548_/Y _06549_/A _06548_/A _06550_/Y vssd1 vssd1 vccd1 vccd1
+ _06555_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09274_ _09276_/C _09274_/B _09274_/C vssd1 vssd1 vccd1 vccd1 _09274_/Y sky130_fd_sc_hd__nor3_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06486_ _06440_/X _06483_/Y _06420_/X _06485_/X vssd1 vssd1 vccd1 vccd1 _13230_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_178_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08225_ _13092_/Q _10433_/B _13087_/Q _10418_/A _08224_/X vssd1 vssd1 vccd1 vccd1
+ _08238_/B sky130_fd_sc_hd__a221o_1
X_08156_ _12822_/Q vssd1 vssd1 vccd1 vccd1 _10454_/B sky130_fd_sc_hd__inv_2
XFILLER_101_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07107_ _07084_/Y _07285_/A _13146_/Q _11514_/X _07106_/X vssd1 vssd1 vccd1 vccd1
+ _13146_/D sky130_fd_sc_hd__a32o_1
XFILLER_106_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08087_ _08284_/A vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07038_ _11970_/X _08562_/B vssd1 vssd1 vccd1 vccd1 _07059_/A sky130_fd_sc_hd__or2_4
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08989_ _12940_/Q vssd1 vssd1 vccd1 vccd1 _08989_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10951_ _10944_/Y _10945_/Y _10895_/Y _10950_/X vssd1 vssd1 vccd1 vccd1 _10977_/D
+ sky130_fd_sc_hd__a31oi_4
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10882_ _12523_/Q _12335_/Q _10873_/Y _10876_/Y vssd1 vssd1 vccd1 vccd1 _10882_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12621_ _13254_/CLK _12945_/Q _08917_/X vssd1 vssd1 vccd1 vccd1 _12621_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_25_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12552_ _13254_/CLK _12552_/D _09066_/X vssd1 vssd1 vccd1 vccd1 _12552_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11503_ _10378_/X _09180_/A _11513_/S vssd1 vssd1 vccd1 vccd1 _11503_/X sky130_fd_sc_hd__mux2_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12483_ _12485_/CLK _12483_/D vssd1 vssd1 vccd1 vccd1 _12483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11434_ _12909_/Q _09179_/B _11443_/S vssd1 vssd1 vccd1 vccd1 _11434_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11365_ _12444_/Q _11364_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _11365_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_4_wb_clk_i _12844_/CLK vssd1 vssd1 vccd1 vccd1 _13081_/CLK sky130_fd_sc_hd__clkbuf_16
X_13104_ _12167_/X _13104_/D _07226_/X vssd1 vssd1 vccd1 vccd1 _13104_/Q sky130_fd_sc_hd__dfrtp_1
X_10316_ _10324_/A vssd1 vssd1 vccd1 vccd1 _10371_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_140_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11296_ vssd1 vssd1 vccd1 vccd1 _11296_/HI _11296_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13035_ _12164_/X _13035_/D _07426_/X vssd1 vssd1 vccd1 vccd1 _13035_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10247_ _13019_/Q _10228_/X _13052_/Q _10229_/X vssd1 vssd1 vccd1 vccd1 _10247_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10178_ _13262_/Q vssd1 vssd1 vccd1 vccd1 _10178_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12819_ _12169_/X _12819_/D _08318_/X vssd1 vssd1 vccd1 vccd1 _12819_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06340_ _06117_/Y _06118_/Y _06122_/Y vssd1 vssd1 vccd1 vccd1 _06340_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06271_ _12045_/S vssd1 vssd1 vccd1 vccd1 _06271_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_147_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08010_ _08018_/A vssd1 vssd1 vccd1 vccd1 _08010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09961_ _08745_/Y _09897_/A _06188_/X _09892_/A _09941_/A vssd1 vssd1 vccd1 vccd1
+ _09961_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_170_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08912_ _08912_/A vssd1 vssd1 vccd1 vccd1 _08912_/X sky130_fd_sc_hd__clkbuf_1
X_09892_ _09892_/A vssd1 vssd1 vccd1 vccd1 _09892_/X sky130_fd_sc_hd__buf_2
XFILLER_97_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08843_ _07746_/X _06283_/Y _08837_/X _12651_/Q vssd1 vssd1 vccd1 vccd1 _12651_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08774_ _12676_/Q vssd1 vssd1 vccd1 vccd1 _08774_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07725_ _12311_/Q vssd1 vssd1 vccd1 vccd1 _07726_/A sky130_fd_sc_hd__inv_2
XFILLER_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07656_ _07659_/A _12953_/Q vssd1 vssd1 vccd1 vccd1 _07657_/D sky130_fd_sc_hd__nand2_1
XPHY_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_74_wb_clk_i _13219_/CLK vssd1 vssd1 vccd1 vccd1 _13205_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06607_ _13218_/Q vssd1 vssd1 vccd1 vccd1 _06607_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07587_ _09271_/A vssd1 vssd1 vccd1 vccd1 _09269_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_179_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09326_ _12363_/Q vssd1 vssd1 vccd1 vccd1 _09327_/B sky130_fd_sc_hd__inv_2
XFILLER_167_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06538_ _13254_/Q _11083_/A _06427_/X _06982_/A _06537_/Y vssd1 vssd1 vccd1 vccd1
+ _11135_/A sky130_fd_sc_hd__o221a_2
XFILLER_139_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09257_ _12452_/Q _09250_/X _09243_/D _09251_/X vssd1 vssd1 vccd1 vccd1 _12452_/D
+ sky130_fd_sc_hd__a22o_1
X_06469_ _06917_/A vssd1 vssd1 vccd1 vccd1 _11107_/A sky130_fd_sc_hd__inv_2
XFILLER_166_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08208_ _08197_/Y _08113_/X _13105_/Q _10467_/A _08207_/X vssd1 vssd1 vccd1 vccd1
+ _08208_/X sky130_fd_sc_hd__o221a_1
XFILLER_138_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09188_ _10796_/D vssd1 vssd1 vccd1 vccd1 _11817_/S sky130_fd_sc_hd__clkinv_16
XFILLER_107_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08139_ _13134_/Q _10460_/A _13129_/Q _10444_/A vssd1 vssd1 vccd1 vccd1 _08139_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11150_ vssd1 vssd1 vccd1 vccd1 _11150_/HI _11150_/LO sky130_fd_sc_hd__conb_1
XFILLER_135_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10101_ _12848_/Q vssd1 vssd1 vccd1 vccd1 _10101_/Y sky130_fd_sc_hd__inv_2
X_11081_ _10763_/X _11071_/X _06379_/X _11058_/X _11072_/X vssd1 vssd1 vccd1 vccd1
+ _11081_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput201 la_oenb[15] vssd1 vssd1 vccd1 vccd1 input201/X sky130_fd_sc_hd__buf_1
XFILLER_103_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput212 la_oenb[25] vssd1 vssd1 vccd1 vccd1 input212/X sky130_fd_sc_hd__buf_1
X_10032_ _10032_/A vssd1 vssd1 vccd1 vccd1 _10032_/X sky130_fd_sc_hd__buf_2
Xinput223 la_oenb[35] vssd1 vssd1 vccd1 vccd1 input223/X sky130_fd_sc_hd__buf_1
Xinput234 la_oenb[45] vssd1 vssd1 vccd1 vccd1 input234/X sky130_fd_sc_hd__buf_1
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput245 la_oenb[55] vssd1 vssd1 vccd1 vccd1 input245/X sky130_fd_sc_hd__buf_1
XFILLER_49_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput256 la_oenb[65] vssd1 vssd1 vccd1 vccd1 input256/X sky130_fd_sc_hd__buf_1
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput267 la_oenb[75] vssd1 vssd1 vccd1 vccd1 input267/X sky130_fd_sc_hd__buf_1
Xinput278 la_oenb[85] vssd1 vssd1 vccd1 vccd1 input278/X sky130_fd_sc_hd__buf_1
XFILLER_5_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput289 la_oenb[95] vssd1 vssd1 vccd1 vccd1 input289/X sky130_fd_sc_hd__buf_1
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11983_ _12615_/Q _09259_/Y _12607_/Q vssd1 vssd1 vccd1 vccd1 _11983_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _12468_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10934_ _10934_/A vssd1 vssd1 vccd1 vccd1 _10947_/B sky130_fd_sc_hd__inv_2
XFILLER_44_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10865_ _10854_/Y _10855_/Y _10849_/Y _10850_/Y vssd1 vssd1 vccd1 vccd1 _10865_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_25_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12604_ _12974_/CLK _12604_/D vssd1 vssd1 vccd1 vccd1 _12604_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _10796_/A _10796_/B _10796_/C _10796_/D vssd1 vssd1 vccd1 vccd1 _12548_/D
+ sky130_fd_sc_hd__nor4_2
XFILLER_157_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _12535_/CLK _12535_/D vssd1 vssd1 vccd1 vccd1 _12535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12466_ _12985_/CLK _12466_/D vssd1 vssd1 vccd1 vccd1 _12466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ _10315_/X _09184_/B _11417_/S vssd1 vssd1 vccd1 vccd1 _11417_/X sky130_fd_sc_hd__mux2_1
X_12397_ _12415_/CLK _12397_/D vssd1 vssd1 vccd1 vccd1 _12397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11348_ _11878_/S _09296_/X _11348_/S vssd1 vssd1 vccd1 vccd1 _11348_/X sky130_fd_sc_hd__mux2_2
XFILLER_126_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11279_ vssd1 vssd1 vccd1 vccd1 _11279_/HI _11279_/LO sky130_fd_sc_hd__conb_1
X_13018_ _12164_/X _13018_/D _07469_/X vssd1 vssd1 vccd1 vccd1 _13018_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07510_ _07609_/A _07510_/B vssd1 vssd1 vccd1 vccd1 _13006_/D sky130_fd_sc_hd__nor2_1
X_08490_ _08441_/Y _10397_/A _08488_/Y _12915_/Q _08489_/X vssd1 vssd1 vccd1 vccd1
+ _08493_/C sky130_fd_sc_hd__o221a_1
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07441_ _07443_/A vssd1 vssd1 vccd1 vccd1 _07441_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07372_ _11430_/X _07368_/X _13054_/Q _07369_/X vssd1 vssd1 vccd1 vccd1 _13054_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09111_ _12527_/Q _09107_/X input337/X _09108_/X vssd1 vssd1 vccd1 vccd1 _12527_/D
+ sky130_fd_sc_hd__a22o_1
X_06323_ _06323_/A vssd1 vssd1 vccd1 vccd1 _06323_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_149_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09042_ _09071_/B _09042_/B _09072_/C vssd1 vssd1 vccd1 vccd1 _09433_/B sky130_fd_sc_hd__or3_4
X_06254_ _12735_/Q _12703_/Q _06259_/A _06253_/Y vssd1 vssd1 vccd1 vccd1 _06254_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06185_ _06185_/A _06209_/A _06197_/B vssd1 vssd1 vccd1 vccd1 _06185_/X sky130_fd_sc_hd__or3_1
XFILLER_117_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ _08794_/Y _09943_/X _06265_/X _09938_/X _09941_/X vssd1 vssd1 vccd1 vccd1
+ _09944_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_132_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09875_ _09873_/Y _09874_/X _09873_/Y _09874_/X vssd1 vssd1 vccd1 vccd1 _09879_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08826_ _08836_/A vssd1 vssd1 vccd1 vccd1 _08826_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _08756_/Y _08565_/X _06204_/X _08742_/X vssd1 vssd1 vccd1 vccd1 _12681_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _12957_/Q _07707_/X _12956_/Q _07705_/X _07703_/X vssd1 vssd1 vccd1 vccd1
+ _12957_/D sky130_fd_sc_hd__o221a_1
XPHY_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08699_/A sky130_fd_sc_hd__buf_2
XFILLER_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ _12955_/Q vssd1 vssd1 vccd1 vccd1 _07665_/A sky130_fd_sc_hd__inv_2
XPHY_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10650_ _12424_/Q vssd1 vssd1 vccd1 vccd1 _10650_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09309_ _09030_/A _09288_/Y _07702_/A _09278_/Y _09292_/B vssd1 vssd1 vccd1 vccd1
+ _12309_/D sky130_fd_sc_hd__o221ai_1
XFILLER_22_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10581_ _10583_/A _11388_/X vssd1 vssd1 vccd1 vccd1 _10581_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_167_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12320_ _12987_/CLK _12320_/D vssd1 vssd1 vccd1 vccd1 _12320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12251_ _12780_/Q _12853_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12251_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11202_ vssd1 vssd1 vccd1 vccd1 _11202_/HI _11202_/LO sky130_fd_sc_hd__conb_1
XFILLER_119_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12182_ _12756_/Q _10688_/X _12755_/Q vssd1 vssd1 vccd1 vccd1 _12182_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11133_ _10758_/X _11100_/X _13249_/Q _11107_/X _11108_/X vssd1 vssd1 vccd1 vccd1
+ _11133_/X sky130_fd_sc_hd__a221o_1
XFILLER_77_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11064_ _10686_/X _10759_/X _06410_/X _10760_/X _10761_/X vssd1 vssd1 vccd1 vccd1
+ _11064_/X sky130_fd_sc_hd__a221o_1
XFILLER_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10015_ _12925_/Q _10015_/B vssd1 vssd1 vccd1 vccd1 _10015_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11966_ _11965_/X _09264_/X _11966_/S vssd1 vssd1 vccd1 vccd1 _11966_/X sky130_fd_sc_hd__mux2_1
X_10917_ _10915_/A _10916_/A _10921_/C _10916_/Y vssd1 vssd1 vccd1 vccd1 _12341_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11897_ _10771_/X _10774_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _11897_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10848_ _10847_/A _10846_/Y _10864_/B _10846_/A vssd1 vssd1 vccd1 vccd1 _12331_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10779_ _10779_/A vssd1 vssd1 vccd1 vccd1 _10779_/X sky130_fd_sc_hd__buf_2
XFILLER_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12518_ _12801_/CLK _12518_/D vssd1 vssd1 vccd1 vccd1 _12518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12449_ _12492_/CLK _12449_/D vssd1 vssd1 vccd1 vccd1 _12449_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_172_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput505 _11254_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__clkbuf_2
Xoutput516 _11264_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput527 _11274_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput538 _11284_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__clkbuf_2
Xoutput549 _11294_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__clkbuf_2
XFILLER_125_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07990_ _07990_/A vssd1 vssd1 vccd1 vccd1 _07990_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_114_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06941_ _06941_/A vssd1 vssd1 vccd1 vccd1 _13182_/D sky130_fd_sc_hd__inv_2
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09660_ _09673_/B _09659_/X _09491_/A vssd1 vssd1 vccd1 vccd1 _09660_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_80_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06872_ _12039_/X _06872_/B vssd1 vssd1 vccd1 vccd1 _06872_/X sky130_fd_sc_hd__or2_1
XFILLER_68_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08611_ _11946_/X _08608_/X _12737_/Q _08610_/X vssd1 vssd1 vccd1 vccd1 _12737_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09591_ _09607_/B vssd1 vssd1 vccd1 vccd1 _09594_/A sky130_fd_sc_hd__inv_2
XFILLER_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08542_ _12754_/Q _08541_/C _08541_/X vssd1 vssd1 vccd1 vccd1 _12754_/D sky130_fd_sc_hd__a21bo_1
XFILLER_36_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08473_ _08468_/X _08473_/B _08473_/C _08473_/D vssd1 vssd1 vccd1 vccd1 _08473_/X
+ sky130_fd_sc_hd__and4b_1
XPHY_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07424_ _07428_/A vssd1 vssd1 vccd1 vccd1 _07424_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07355_ _11437_/X _07353_/X _13061_/Q _07354_/X vssd1 vssd1 vccd1 vccd1 _13061_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06306_ _06306_/A vssd1 vssd1 vccd1 vccd1 _06306_/X sky130_fd_sc_hd__clkbuf_2
X_07286_ _09183_/A vssd1 vssd1 vccd1 vccd1 _09242_/A sky130_fd_sc_hd__buf_6
XFILLER_108_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09025_ _12602_/Q vssd1 vssd1 vccd1 vccd1 _10015_/B sky130_fd_sc_hd__clkbuf_2
X_06237_ _06051_/A _06184_/X _06051_/A _06184_/X vssd1 vssd1 vccd1 vccd1 _06237_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_85_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06168_ _08996_/D vssd1 vssd1 vccd1 vccd1 _06214_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06099_ _12725_/Q vssd1 vssd1 vccd1 vccd1 _06099_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _09925_/Y _09922_/X _06295_/A _09915_/X _09926_/X vssd1 vssd1 vccd1 vccd1
+ _09927_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09858_ _13234_/Q _09857_/B _09857_/Y vssd1 vssd1 vccd1 vccd1 _09866_/B sky130_fd_sc_hd__o21ai_2
XFILLER_105_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08809_ _08839_/A vssd1 vssd1 vccd1 vccd1 _08823_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09789_ _06577_/Y _09788_/X _06577_/Y _09788_/X vssd1 vssd1 vccd1 vccd1 _09790_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _09889_/X _12845_/Q _11831_/S vssd1 vssd1 vccd1 vccd1 _11820_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11751_ _11376_/X _12472_/Q _12103_/S vssd1 vssd1 vccd1 vccd1 _11751_/X sky130_fd_sc_hd__mux2_1
XPHY_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10702_ _06410_/X _11058_/A _10686_/X _11071_/A _06637_/Y vssd1 vssd1 vccd1 vccd1
+ _10702_/X sky130_fd_sc_hd__o221a_1
XPHY_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11682_ _11681_/X _11378_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12383_/D sky130_fd_sc_hd__mux2_1
XPHY_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _08926_/A _08926_/B _08927_/B vssd1 vssd1 vccd1 vccd1 _10633_/X sky130_fd_sc_hd__a21bo_1
XFILLER_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10564_ _10564_/A vssd1 vssd1 vccd1 vccd1 _11390_/S sky130_fd_sc_hd__inv_2
XFILLER_154_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12303_ _12977_/CLK _12303_/D vssd1 vssd1 vccd1 vccd1 _12303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13283_ _13283_/CLK _13283_/D _06194_/X vssd1 vssd1 vccd1 vccd1 _13283_/Q sky130_fd_sc_hd__dfrtp_1
X_10495_ _12500_/Q _09139_/B _09140_/B vssd1 vssd1 vccd1 vccd1 _10495_/X sky130_fd_sc_hd__a21bo_1
XFILLER_6_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12234_ _12233_/X _12637_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__mux2_2
XFILLER_182_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12165_ _12165_/A0 input23/X _12843_/Q vssd1 vssd1 vccd1 vccd1 _12165_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11116_ _10755_/A _11054_/A _13250_/Q _11055_/A _11899_/X vssd1 vssd1 vccd1 vccd1
+ _11116_/X sky130_fd_sc_hd__a221o_1
XFILLER_2_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12096_ _12095_/X _12448_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11047_ _11033_/X _11037_/X _06397_/X _07020_/X _11038_/X vssd1 vssd1 vccd1 vccd1
+ _11047_/X sky130_fd_sc_hd__a221o_1
XFILLER_65_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 io_in[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XFILLER_92_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12998_ _13001_/CLK _12998_/D vssd1 vssd1 vccd1 vccd1 _12998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11949_ _09796_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11949_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07140_ _07152_/A vssd1 vssd1 vccd1 vccd1 _07140_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07071_ _07078_/A vssd1 vssd1 vccd1 vccd1 _07071_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06022_ _06281_/A vssd1 vssd1 vccd1 vccd1 _06022_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput368 _12964_/Q vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__clkbuf_2
Xoutput379 _11164_/LO vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07973_ _07976_/A vssd1 vssd1 vccd1 vccd1 _07996_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09712_ _09711_/A _09711_/B _09711_/Y vssd1 vssd1 vccd1 vccd1 _09747_/A sky130_fd_sc_hd__a21oi_4
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06924_ _11995_/X _06924_/B vssd1 vssd1 vccd1 vccd1 _06924_/X sky130_fd_sc_hd__or2_2
XFILLER_56_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09643_ _09643_/A _09643_/B vssd1 vssd1 vccd1 vccd1 _09659_/A sky130_fd_sc_hd__nor2_2
XFILLER_110_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06855_ _12027_/X _06819_/X _12027_/X _06819_/X vssd1 vssd1 vccd1 vccd1 _06864_/B
+ sky130_fd_sc_hd__a2bb2oi_4
XFILLER_28_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09574_ _09574_/A _09574_/B _09530_/A vssd1 vssd1 vccd1 vccd1 _09574_/X sky130_fd_sc_hd__or3b_1
X_06786_ _12016_/X _12012_/X _06785_/X vssd1 vssd1 vccd1 vccd1 _06786_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08525_ _08519_/X _12244_/X _08514_/X _12759_/Q vssd1 vssd1 vccd1 vccd1 _12759_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08456_ _08445_/Y _07800_/X _13065_/Q _10380_/A _08455_/X vssd1 vssd1 vccd1 vccd1
+ _08456_/X sky130_fd_sc_hd__o221a_1
XPHY_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07407_ _07403_/Y _08251_/A _13146_/Q _11417_/X _07406_/X vssd1 vssd1 vccd1 vccd1
+ _13041_/D sky130_fd_sc_hd__a32o_1
XFILLER_17_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08387_ _08657_/A vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__buf_2
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07338_ _07368_/A vssd1 vssd1 vccd1 vccd1 _07338_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07269_ _07362_/A vssd1 vssd1 vccd1 vccd1 _07280_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ _09008_/A _09008_/B _11644_/X vssd1 vssd1 vccd1 vccd1 _12588_/D sky130_fd_sc_hd__and3_1
XFILLER_152_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10280_ _13268_/Q vssd1 vssd1 vccd1 vccd1 _10280_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _12166_/X _12921_/D _07899_/X vssd1 vssd1 vccd1 vccd1 _12921_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12852_/CLK _12852_/D _08088_/X vssd1 vssd1 vccd1 vccd1 _12852_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _10679_/X _10792_/B _11803_/S vssd1 vssd1 vccd1 vccd1 _11803_/X sky130_fd_sc_hd__mux2_1
XPHY_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12942_/CLK _12783_/D _08412_/X vssd1 vssd1 vccd1 vccd1 _12783_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11734_ _11733_/X _11414_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12443_/D sky130_fd_sc_hd__mux2_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11665_ _11381_/X _09185_/C _11675_/S vssd1 vssd1 vccd1 vccd1 _11665_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10616_ _12411_/D _10617_/A vssd1 vssd1 vccd1 vccd1 _10616_/Y sky130_fd_sc_hd__nor2_1
XPHY_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11596_ _10452_/Y _09179_/A _11603_/S vssd1 vssd1 vccd1 vccd1 _11596_/X sky130_fd_sc_hd__mux2_1
XPHY_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10547_ _11358_/X _10554_/B vssd1 vssd1 vccd1 vccd1 _10547_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13266_ _13269_/CLK _13266_/D _06293_/X vssd1 vssd1 vccd1 vccd1 _13266_/Q sky130_fd_sc_hd__dfrtp_1
X_10478_ _10480_/B vssd1 vssd1 vccd1 vccd1 _10478_/Y sky130_fd_sc_hd__inv_2
X_12217_ _06316_/X _13154_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12217_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13197_ _13201_/CLK _13197_/D _06803_/X vssd1 vssd1 vccd1 vccd1 _13197_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12148_ _09997_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12148_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12079_ _12078_/X _12446_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12079_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06640_ _11901_/X _12196_/X _06639_/X vssd1 vssd1 vccd1 vccd1 _06640_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06571_ _12179_/X _06543_/X _12179_/X _06543_/X vssd1 vssd1 vccd1 vccd1 _06576_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_17_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08310_ _12823_/Q _11598_/X _08321_/S vssd1 vssd1 vccd1 vccd1 _12823_/D sky130_fd_sc_hd__mux2_1
X_09290_ _09269_/A _08984_/Y _13006_/Q _09288_/B _09027_/B vssd1 vssd1 vccd1 vccd1
+ _09290_/X sky130_fd_sc_hd__o32a_1
XFILLER_166_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ _13111_/Q _10482_/A _13106_/Q _08164_/Y vssd1 vssd1 vccd1 vccd1 _08246_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_177_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08172_ _13130_/Q _10449_/B _13133_/Q _10454_/A _08171_/X vssd1 vssd1 vccd1 vccd1
+ _08175_/C sky130_fd_sc_hd__o221a_1
XFILLER_118_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07123_ _11543_/X _07113_/X _13142_/Q _07116_/X vssd1 vssd1 vccd1 vccd1 _13142_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07054_ _07053_/X _07040_/X _06295_/Y _13158_/Q _07042_/X vssd1 vssd1 vccd1 vccd1
+ _13158_/D sky130_fd_sc_hd__a32o_1
XFILLER_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06005_ _13286_/Q vssd1 vssd1 vccd1 vccd1 _06005_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_28_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12430_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_173_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07956_ _12898_/Q _11487_/X _07962_/S vssd1 vssd1 vccd1 vccd1 _12898_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06907_ _06907_/A vssd1 vssd1 vccd1 vccd1 _13186_/D sky130_fd_sc_hd__inv_2
XFILLER_96_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07887_ _07886_/Y input1/X _07886_/Y input1/X vssd1 vssd1 vccd1 vccd1 _07887_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09626_ _13159_/Q vssd1 vssd1 vccd1 vccd1 _09626_/Y sky130_fd_sc_hd__inv_2
X_06838_ _06435_/X _12189_/X _06436_/X _13194_/Q vssd1 vssd1 vccd1 vccd1 _13194_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_56_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09557_ _09522_/A _09574_/A _09522_/B _09574_/A _09556_/Y vssd1 vssd1 vccd1 vccd1
+ _09558_/B sky130_fd_sc_hd__o221a_1
XFILLER_110_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06769_ _06769_/A vssd1 vssd1 vccd1 vccd1 _06769_/X sky130_fd_sc_hd__clkbuf_4
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08508_ _08504_/X _12258_/X _08499_/X _12766_/Q vssd1 vssd1 vccd1 vccd1 _12766_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_169_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09488_ _13167_/Q _13166_/Q _13167_/Q _13166_/Q vssd1 vssd1 vccd1 vccd1 _09488_/X
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08439_ _12772_/Q _08417_/A _07568_/X _08418_/A vssd1 vssd1 vccd1 vccd1 _12772_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11450_ _12893_/Q _09184_/A _11459_/S vssd1 vssd1 vccd1 vccd1 _11450_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10401_ input23/X vssd1 vssd1 vccd1 vccd1 _10401_/Y sky130_fd_sc_hd__inv_2
X_11381_ _10568_/X _12397_/D _11392_/S vssd1 vssd1 vccd1 vccd1 _11381_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _12168_/X _13120_/D _07179_/X vssd1 vssd1 vccd1 vccd1 _13120_/Q sky130_fd_sc_hd__dfrtp_2
X_10332_ _12898_/Q _10329_/Y _10333_/B _10320_/X vssd1 vssd1 vccd1 vccd1 _10332_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13051_ _12165_/X _13051_/D _07379_/X vssd1 vssd1 vccd1 vccd1 _13051_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ _13267_/Q vssd1 vssd1 vccd1 vccd1 _10263_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12002_ _11105_/X _11097_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _12002_/X sky130_fd_sc_hd__mux2_2
XFILLER_106_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10194_ _07803_/Y _10151_/X _10193_/X vssd1 vssd1 vccd1 vccd1 _10194_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_94_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12904_ _12166_/X _12904_/D _07939_/X vssd1 vssd1 vccd1 vccd1 _12904_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ _12169_/X _12835_/D _08268_/X vssd1 vssd1 vccd1 vccd1 _12835_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12766_ _12769_/CLK _12766_/D _08507_/X vssd1 vssd1 vccd1 vccd1 _12766_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11717_ _10648_/Y _10649_/Y _11818_/S vssd1 vssd1 vccd1 vccd1 _11717_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12697_ _12719_/CLK _12697_/D _08710_/X vssd1 vssd1 vccd1 vccd1 _12697_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _10518_/X _12933_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11648_/X sky130_fd_sc_hd__mux2_1
Xinput12 io_in[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_4
Xinput23 io_in[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_4
XFILLER_168_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput34 io_in[5] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_1
XFILLER_156_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput45 la_data_in[105] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_1
XFILLER_190_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11579_ _10404_/Y _09184_/A _11592_/S vssd1 vssd1 vccd1 vccd1 _11579_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput56 la_data_in[115] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_1
XFILLER_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput67 la_data_in[125] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_1
Xinput78 la_data_in[1] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__buf_4
XFILLER_122_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput89 la_data_in[2] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__buf_1
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13249_ _13249_/CLK _13249_/D _06374_/X vssd1 vssd1 vccd1 vccd1 _13249_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07810_ _12906_/Q vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__inv_2
XFILLER_85_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08790_ _12671_/Q vssd1 vssd1 vccd1 vccd1 _08790_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater613 _11603_/S vssd1 vssd1 vccd1 vccd1 _11592_/S sky130_fd_sc_hd__buf_4
Xrepeater624 _11422_/S vssd1 vssd1 vccd1 vccd1 _11449_/S sky130_fd_sc_hd__clkbuf_4
Xrepeater635 input356/X vssd1 vssd1 vccd1 vccd1 _09185_/B sky130_fd_sc_hd__buf_8
X_07741_ _12615_/Q vssd1 vssd1 vccd1 vccd1 _08837_/A sky130_fd_sc_hd__buf_2
XFILLER_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater646 _07975_/A vssd1 vssd1 vccd1 vccd1 _10528_/B sky130_fd_sc_hd__buf_8
XFILLER_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07672_ _07685_/C _07676_/A _07672_/C _07689_/D vssd1 vssd1 vccd1 vccd1 _07679_/A
+ sky130_fd_sc_hd__or4b_4
Xclkbuf_leaf_146_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12875_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09411_ _12396_/D vssd1 vssd1 vccd1 vccd1 _09411_/Y sky130_fd_sc_hd__inv_2
X_06623_ _06435_/X _12191_/X _06436_/X _13217_/Q vssd1 vssd1 vccd1 vccd1 _13217_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09342_ _12402_/Q vssd1 vssd1 vccd1 vccd1 _09342_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06554_ _06580_/A vssd1 vssd1 vccd1 vccd1 _06554_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09273_ _12299_/Q _12304_/Q _12300_/Q _12301_/Q vssd1 vssd1 vccd1 vccd1 _09274_/C
+ sky130_fd_sc_hd__or4_4
X_06485_ _12044_/X _12043_/X _12041_/X _06484_/X vssd1 vssd1 vccd1 vccd1 _06485_/X
+ sky130_fd_sc_hd__o22a_1
X_08224_ _13102_/Q _10460_/A _13097_/Q _10444_/A vssd1 vssd1 vccd1 vccd1 _08224_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08155_ _08141_/Y _10405_/A _13139_/Q _08154_/Y vssd1 vssd1 vccd1 vccd1 _08162_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07106_ _13079_/Q _07284_/A vssd1 vssd1 vccd1 vccd1 _07106_/X sky130_fd_sc_hd__or2_1
XFILLER_161_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08086_ _12853_/Q _08082_/X _07287_/X _08083_/X vssd1 vssd1 vccd1 vccd1 _12853_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_161_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07037_ _07069_/A vssd1 vssd1 vccd1 vccd1 _07037_/X sky130_fd_sc_hd__buf_2
XFILLER_161_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08988_ _12964_/Q _12963_/Q _08995_/C vssd1 vssd1 vccd1 vccd1 _08988_/X sky130_fd_sc_hd__and3_1
XFILLER_57_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07939_ _07945_/A vssd1 vssd1 vccd1 vccd1 _07939_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10950_ _12533_/Q _12345_/Q _10949_/X vssd1 vssd1 vccd1 vccd1 _10950_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ _09609_/A _09632_/A vssd1 vssd1 vccd1 vccd1 _09609_/X sky130_fd_sc_hd__or2_1
X_10881_ _10879_/Y _10880_/Y _12524_/Q _12336_/Q vssd1 vssd1 vccd1 vccd1 _10888_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _12620_/CLK _12620_/D vssd1 vssd1 vccd1 vccd1 _12620_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _12169_/A0 _12551_/D _09067_/X vssd1 vssd1 vccd1 vccd1 _12551_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11502_ _10374_/X _09180_/B _11513_/S vssd1 vssd1 vccd1 vccd1 _11502_/X sky130_fd_sc_hd__mux2_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12482_ _12485_/CLK _12482_/D vssd1 vssd1 vccd1 vccd1 _12482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11433_ _12908_/Q _10528_/B _11433_/S vssd1 vssd1 vccd1 vccd1 _11433_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11364_ _11363_/X _12444_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _11364_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10315_ _13146_/Q _12551_/Q vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__or2_1
X_13103_ _12167_/X _13103_/D _07228_/X vssd1 vssd1 vccd1 vccd1 _13103_/Q sky130_fd_sc_hd__dfrtp_1
X_11295_ vssd1 vssd1 vccd1 vccd1 _11295_/HI _11295_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13034_ _12164_/X _13034_/D _07428_/X vssd1 vssd1 vccd1 vccd1 _13034_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10246_ _13092_/Q _10228_/X _13124_/Q _10229_/X vssd1 vssd1 vccd1 vccd1 _10246_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10177_ _12661_/Q vssd1 vssd1 vccd1 vccd1 _10177_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12818_ _12169_/X _12818_/D _08320_/X vssd1 vssd1 vccd1 vccd1 _12818_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12749_ _12749_/CLK _12749_/D _08569_/X vssd1 vssd1 vccd1 vccd1 _12749_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06270_ _06064_/A _06064_/B _06134_/A _06134_/Y _06069_/A vssd1 vssd1 vccd1 vccd1
+ _12045_/S sky130_fd_sc_hd__a32o_2
XFILLER_175_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09960_ _08748_/Y _09897_/A _06192_/X _09892_/A _09941_/A vssd1 vssd1 vccd1 vccd1
+ _09960_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08911_ _08898_/X _06342_/Y _08908_/X _12624_/Q vssd1 vssd1 vccd1 vccd1 _12624_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_103_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09891_ _09891_/A vssd1 vssd1 vccd1 vccd1 _09892_/A sky130_fd_sc_hd__buf_2
XFILLER_97_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08842_ _08851_/A vssd1 vssd1 vccd1 vccd1 _08842_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08773_ _08789_/A vssd1 vssd1 vccd1 vccd1 _08773_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07724_ _07678_/A _07717_/X _12946_/Q _07693_/X _09288_/A vssd1 vssd1 vccd1 vccd1
+ _12947_/D sky130_fd_sc_hd__o221a_1
XFILLER_26_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07655_ _07642_/B _07646_/D _12957_/Q _07665_/A vssd1 vssd1 vccd1 vccd1 _07684_/A
+ sky130_fd_sc_hd__and4bb_1
XPHY_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06606_ _06650_/A vssd1 vssd1 vccd1 vccd1 _06606_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07586_ _12602_/Q vssd1 vssd1 vccd1 vccd1 _09271_/A sky130_fd_sc_hd__inv_2
XFILLER_129_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09325_ _12364_/Q vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__inv_2
XFILLER_179_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06537_ _12089_/X vssd1 vssd1 vccd1 vccd1 _06537_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09256_ _12453_/Q _09250_/X _09243_/C _09251_/X vssd1 vssd1 vccd1 vccd1 _12453_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06468_ _06468_/A _12766_/Q vssd1 vssd1 vccd1 vccd1 _06917_/A sky130_fd_sc_hd__or2b_2
XFILLER_193_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08207_ _08205_/Y _08128_/X _08206_/Y _12813_/Q vssd1 vssd1 vccd1 vccd1 _08207_/X
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_43_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12984_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09187_ _09187_/A _09187_/B _09187_/C _10535_/A vssd1 vssd1 vccd1 vccd1 _10796_/D
+ sky130_fd_sc_hd__or4_4
X_06399_ _06412_/A vssd1 vssd1 vccd1 vccd1 _06399_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08138_ _12819_/Q vssd1 vssd1 vccd1 vccd1 _10444_/A sky130_fd_sc_hd__inv_2
XFILLER_119_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08069_ _12860_/Q _08066_/X _07975_/X _08068_/X vssd1 vssd1 vccd1 vccd1 _12860_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_161_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10100_ _10098_/Y _10023_/X _10099_/Y _10025_/X vssd1 vssd1 vccd1 vccd1 _10107_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11080_ _06371_/X _11045_/X _08535_/A _10755_/X _07030_/X vssd1 vssd1 vccd1 vccd1
+ _11080_/X sky130_fd_sc_hd__a32o_1
XFILLER_1_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput202 la_oenb[16] vssd1 vssd1 vccd1 vccd1 input202/X sky130_fd_sc_hd__buf_1
XFILLER_1_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10031_ _13255_/Q vssd1 vssd1 vccd1 vccd1 _10031_/Y sky130_fd_sc_hd__inv_2
Xinput213 la_oenb[26] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__buf_1
XFILLER_102_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput224 la_oenb[36] vssd1 vssd1 vccd1 vccd1 input224/X sky130_fd_sc_hd__buf_1
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput235 la_oenb[46] vssd1 vssd1 vccd1 vccd1 input235/X sky130_fd_sc_hd__buf_1
XFILLER_124_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput246 la_oenb[56] vssd1 vssd1 vccd1 vccd1 input246/X sky130_fd_sc_hd__buf_1
XFILLER_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput257 la_oenb[66] vssd1 vssd1 vccd1 vccd1 input257/X sky130_fd_sc_hd__buf_1
XFILLER_5_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput268 la_oenb[76] vssd1 vssd1 vccd1 vccd1 input268/X sky130_fd_sc_hd__buf_1
Xinput279 la_oenb[86] vssd1 vssd1 vccd1 vccd1 input279/X sky130_fd_sc_hd__buf_1
XFILLER_91_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11982_ _09037_/X _07520_/Y _11982_/S vssd1 vssd1 vccd1 vccd1 _11982_/X sky130_fd_sc_hd__mux2_4
XFILLER_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10933_ _10933_/A vssd1 vssd1 vccd1 vccd1 _10933_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10864_ _10864_/A _10864_/B _10864_/C _10851_/X vssd1 vssd1 vccd1 vccd1 _10864_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12603_ _13001_/CLK _12603_/D vssd1 vssd1 vccd1 vccd1 _12603_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _12943_/Q _12941_/Q _10795_/C _10795_/D vssd1 vssd1 vccd1 vccd1 _10796_/C
+ sky130_fd_sc_hd__or4_4
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12535_/CLK _12534_/D vssd1 vssd1 vccd1 vccd1 _12534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12465_ _13008_/CLK _12465_/D vssd1 vssd1 vccd1 vccd1 _12465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11416_ _10243_/Y _12798_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11416_/X sky130_fd_sc_hd__mux2_1
X_12396_ _12415_/CLK _12396_/D vssd1 vssd1 vccd1 vccd1 _12396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11347_ input78/X vssd1 vssd1 vccd1 vccd1 _11347_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_153_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11278_ vssd1 vssd1 vccd1 vccd1 _11278_/HI _11278_/LO sky130_fd_sc_hd__conb_1
X_13017_ _12164_/X _13017_/D _07471_/X vssd1 vssd1 vccd1 vccd1 _13017_/Q sky130_fd_sc_hd__dfrtp_1
X_10229_ _10277_/A vssd1 vssd1 vccd1 vccd1 _10229_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07440_ _11471_/X _07429_/X _13030_/Q _07430_/X vssd1 vssd1 vccd1 vccd1 _13030_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07371_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07371_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_188_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09110_ _12528_/Q _09107_/X input338/X _09108_/X vssd1 vssd1 vccd1 vccd1 _12528_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06322_ _06108_/A _06321_/X _06108_/A _06321_/X vssd1 vssd1 vccd1 vccd1 _06323_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_200_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09041_ _09041_/A _09041_/B _07095_/B vssd1 vssd1 vccd1 vccd1 _09072_/C sky130_fd_sc_hd__or3b_1
X_06253_ _06253_/A vssd1 vssd1 vccd1 vccd1 _06253_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06184_ _06209_/C _06173_/X _06181_/X _06182_/X _06183_/X vssd1 vssd1 vccd1 vccd1
+ _06184_/X sky130_fd_sc_hd__o221a_1
XFILLER_171_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09943_ _09952_/A vssd1 vssd1 vccd1 vccd1 _09943_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_161_wb_clk_i clkbuf_opt_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _12541_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09874_ _09862_/Y _06441_/Y _09686_/X _09864_/Y vssd1 vssd1 vccd1 vccd1 _09874_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08825_ _08839_/A vssd1 vssd1 vccd1 vccd1 _08836_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08756_ _12681_/Q vssd1 vssd1 vccd1 vccd1 _08756_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _07717_/A vssd1 vssd1 vccd1 vccd1 _07707_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08687_ _11841_/X _08685_/X _12707_/Q _08686_/X vssd1 vssd1 vccd1 vccd1 _12707_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _07678_/A _07678_/B _07631_/Y _07637_/Y vssd1 vssd1 vccd1 vccd1 _07685_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07569_ _07775_/A vssd1 vssd1 vccd1 vccd1 _07569_/X sky130_fd_sc_hd__buf_2
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09308_ _07719_/A _09278_/Y _09286_/B vssd1 vssd1 vccd1 vccd1 _12310_/D sky130_fd_sc_hd__o21ai_1
XFILLER_167_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10580_ _12401_/D _10578_/Y _10579_/X vssd1 vssd1 vccd1 vccd1 _10580_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09239_ _12461_/Q _09233_/A _07564_/X _09083_/X vssd1 vssd1 vccd1 vccd1 _12461_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_127_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12250_ _12249_/X _12645_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12250_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11201_ vssd1 vssd1 vccd1 vccd1 _11201_/HI _11201_/LO sky130_fd_sc_hd__conb_1
XFILLER_163_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12181_ _10694_/X _10689_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _12181_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11132_ _10742_/A _10759_/A _13251_/Q _11086_/A _12195_/X vssd1 vssd1 vccd1 vccd1
+ _11132_/X sky130_fd_sc_hd__a221o_1
XFILLER_123_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11063_ _10696_/X _10750_/X _06404_/X _10751_/X _10752_/X vssd1 vssd1 vccd1 vccd1
+ _11063_/X sky130_fd_sc_hd__a221o_1
XFILLER_153_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10014_ _12303_/Q _12301_/Q vssd1 vssd1 vccd1 vccd1 _12180_/S sky130_fd_sc_hd__nor2_1
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11965_ _12943_/Q _11964_/X _11969_/S vssd1 vssd1 vccd1 vccd1 _11965_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _10916_/A vssd1 vssd1 vccd1 vccd1 _10916_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11896_ _10782_/Y _10781_/Y _12193_/S vssd1 vssd1 vccd1 vccd1 _11896_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10847_ _10847_/A vssd1 vssd1 vccd1 vccd1 _10864_/B sky130_fd_sc_hd__inv_2
XFILLER_73_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10778_ _10773_/X _10731_/X _06386_/X _10732_/X _10733_/X vssd1 vssd1 vccd1 vccd1
+ _10778_/X sky130_fd_sc_hd__a221o_1
XFILLER_200_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12517_ _12517_/CLK _12517_/D vssd1 vssd1 vccd1 vccd1 _12517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12448_ _12619_/CLK _12448_/D vssd1 vssd1 vccd1 vccd1 _12448_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_201_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput506 _11255_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__clkbuf_2
Xoutput517 _11265_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput528 _11275_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12379_ _12577_/CLK _12379_/D vssd1 vssd1 vccd1 vccd1 _12401_/D sky130_fd_sc_hd__dfxtp_1
Xoutput539 _11285_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__clkbuf_2
XFILLER_119_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06940_ _06841_/A _06935_/B _06938_/Y _06630_/X _09576_/A vssd1 vssd1 vccd1 vccd1
+ _06941_/A sky130_fd_sc_hd__o32a_1
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06871_ _12036_/X vssd1 vssd1 vccd1 vccd1 _06872_/B sky130_fd_sc_hd__inv_2
XFILLER_41_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08610_ _08686_/A vssd1 vssd1 vccd1 vccd1 _08610_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09590_ _09576_/A _09576_/B _09589_/A _09576_/Y _09589_/Y vssd1 vssd1 vccd1 vccd1
+ _09607_/B sky130_fd_sc_hd__o32a_1
XFILLER_48_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08541_ _08849_/A _12045_/X _08541_/C vssd1 vssd1 vccd1 vccd1 _08541_/X sky130_fd_sc_hd__or3_2
XFILLER_78_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08472_ _13053_/Q _10346_/A _08471_/Y _07821_/X vssd1 vssd1 vccd1 vccd1 _08473_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07423_ _11478_/X _07412_/X _13037_/Q _07415_/X vssd1 vssd1 vccd1 vccd1 _13037_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07354_ _07369_/A vssd1 vssd1 vccd1 vccd1 _07354_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06305_ _06305_/A vssd1 vssd1 vccd1 vccd1 _06305_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_176_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07285_ _07285_/A vssd1 vssd1 vccd1 vccd1 _07285_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09024_ _12975_/Q _12974_/Q _12976_/Q vssd1 vssd1 vccd1 vccd1 _09288_/B sky130_fd_sc_hd__nor3_4
X_06236_ _13276_/Q vssd1 vssd1 vccd1 vccd1 _06236_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06167_ _08854_/A vssd1 vssd1 vccd1 vccd1 _08996_/D sky130_fd_sc_hd__buf_6
XFILLER_145_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06098_ _06098_/A vssd1 vssd1 vccd1 vccd1 _06103_/A sky130_fd_sc_hd__inv_2
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09926_ _12888_/Q _09935_/B vssd1 vssd1 vccd1 vccd1 _09926_/X sky130_fd_sc_hd__or2_1
XFILLER_120_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09857_ _13234_/Q _09857_/B vssd1 vssd1 vccd1 vccd1 _09857_/Y sky130_fd_sc_hd__nand2_2
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08808_ _08798_/X _08801_/X _06295_/Y _12665_/Q _08567_/X vssd1 vssd1 vccd1 vccd1
+ _12665_/D sky130_fd_sc_hd__a32o_1
XFILLER_46_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09788_ _06581_/Y _09787_/X _06581_/Y _09787_/X vssd1 vssd1 vccd1 vccd1 _09788_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_65_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _12685_/Q vssd1 vssd1 vccd1 vccd1 _08739_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11749_/X _11374_/X _11774_/S vssd1 vssd1 vccd1 vccd1 _12427_/D sky130_fd_sc_hd__mux2_1
XPHY_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _10701_/A _12757_/Q vssd1 vssd1 vccd1 vccd1 _10701_/Y sky130_fd_sc_hd__nor2_2
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11681_ _11378_/X _09243_/C _11691_/S vssd1 vssd1 vccd1 vccd1 _11681_/X sky130_fd_sc_hd__mux2_1
XPHY_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10632_ _11890_/X _10649_/B vssd1 vssd1 vccd1 vccd1 _10632_/Y sky130_fd_sc_hd__nor2_1
XPHY_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10563_ _12395_/D _12398_/D _10562_/B _10570_/A vssd1 vssd1 vccd1 vccd1 _10564_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _12576_/CLK _12302_/D vssd1 vssd1 vccd1 vccd1 _12302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10494_ _12499_/Q _09138_/B _09139_/B vssd1 vssd1 vccd1 vccd1 _10494_/X sky130_fd_sc_hd__a21bo_1
X_13282_ _13283_/CLK _13282_/D _06202_/X vssd1 vssd1 vccd1 vccd1 _13282_/Q sky130_fd_sc_hd__dfrtp_1
X_12233_ _06271_/Y _13162_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12233_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12164_ _12165_/A0 _10401_/Y _12843_/Q vssd1 vssd1 vccd1 vccd1 _12164_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _10736_/A _11071_/X _13252_/Q _11058_/A _11072_/X vssd1 vssd1 vccd1 vccd1
+ _11115_/X sky130_fd_sc_hd__a221o_1
XFILLER_151_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12095_ _12094_/X _12448_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12095_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11046_ _06389_/X _11045_/X _11032_/X _10779_/X _11034_/X vssd1 vssd1 vccd1 vccd1
+ _11046_/X sky130_fd_sc_hd__a32o_1
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12997_ _13001_/CLK _12997_/D vssd1 vssd1 vccd1 vccd1 _12997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11948_ _09786_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11948_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11879_ _11042_/X _11035_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _11879_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07070_ _07069_/X _07058_/X _06327_/Y _13152_/Q _07059_/X vssd1 vssd1 vccd1 vccd1
+ _13152_/D sky130_fd_sc_hd__a32o_1
XFILLER_199_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06021_ _06314_/A vssd1 vssd1 vccd1 vccd1 _06281_/A sky130_fd_sc_hd__buf_2
XFILLER_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput369 _11151_/HI vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07972_ _09982_/D _09981_/C _08399_/B vssd1 vssd1 vccd1 vccd1 _07976_/A sky130_fd_sc_hd__or3_4
XFILLER_45_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09711_ _09711_/A _09711_/B vssd1 vssd1 vccd1 vccd1 _09711_/Y sky130_fd_sc_hd__nor2_4
XFILLER_101_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06923_ _11992_/X vssd1 vssd1 vccd1 vccd1 _06924_/B sky130_fd_sc_hd__inv_2
XFILLER_45_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09642_ _09640_/A _09640_/B _09641_/Y vssd1 vssd1 vccd1 vccd1 _09643_/B sky130_fd_sc_hd__a21o_1
X_06854_ _06847_/X _06851_/X _06857_/A vssd1 vssd1 vccd1 vccd1 _06864_/A sky130_fd_sc_hd__a21oi_4
XFILLER_95_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06785_ _12037_/X _06785_/B vssd1 vssd1 vccd1 vccd1 _06785_/X sky130_fd_sc_hd__or2_1
X_09573_ _09550_/Y _09566_/A _09563_/A vssd1 vssd1 vccd1 vccd1 _09609_/A sky130_fd_sc_hd__o21ai_1
XFILLER_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08524_ _08533_/A vssd1 vssd1 vccd1 vccd1 _08524_/X sky130_fd_sc_hd__clkbuf_1
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08455_ _08453_/Y _07815_/X _08454_/Y _12902_/Q vssd1 vssd1 vccd1 vccd1 _08455_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07406_ _12841_/Q _08250_/A vssd1 vssd1 vccd1 vccd1 _07406_/X sky130_fd_sc_hd__or2_1
XPHY_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08386_ _12792_/Q _08374_/X _07296_/X _08375_/X vssd1 vssd1 vccd1 vccd1 _12792_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_196_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07337_ _07345_/A vssd1 vssd1 vccd1 vccd1 _07337_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07268_ _07477_/A vssd1 vssd1 vccd1 vccd1 _07362_/A sky130_fd_sc_hd__buf_4
XFILLER_192_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09007_ _09008_/A _09008_/B _11645_/X vssd1 vssd1 vccd1 vccd1 _12589_/D sky130_fd_sc_hd__and3_1
X_06219_ _06215_/Y _06216_/X _06217_/X _06218_/X vssd1 vssd1 vccd1 vccd1 _13280_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_192_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07199_ hold1/X _11558_/S vssd1 vssd1 vccd1 vccd1 _07263_/A sky130_fd_sc_hd__or2_1
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09909_ _12660_/Q vssd1 vssd1 vccd1 vccd1 _09909_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12920_ _12166_/X _12920_/D _07901_/X vssd1 vssd1 vccd1 vccd1 _12920_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _12852_/CLK _12851_/D _08090_/X vssd1 vssd1 vccd1 vccd1 _12851_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _11801_/X _12065_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12440_/D sky130_fd_sc_hd__mux2_1
XPHY_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12942_/CLK _12782_/D _08414_/X vssd1 vssd1 vccd1 vccd1 _12782_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11414_/X _11732_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11733_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11663_/X _11383_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12374_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10615_ _10625_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _10617_/A sky130_fd_sc_hd__or2_2
XFILLER_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11595_ _10448_/X _09179_/B _11603_/S vssd1 vssd1 vccd1 vccd1 _11595_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10546_ _11358_/X vssd1 vssd1 vccd1 vccd1 _10546_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13265_ _13269_/CLK _13265_/D _06297_/X vssd1 vssd1 vccd1 vccd1 _13265_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10477_ _10477_/A _10477_/B vssd1 vssd1 vccd1 vccd1 _10480_/B sky130_fd_sc_hd__or2_1
XFILLER_6_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12216_ _12215_/X _12628_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12216_/X sky130_fd_sc_hd__mux2_1
X_13196_ _13196_/CLK _13196_/D _06806_/X vssd1 vssd1 vccd1 vccd1 _13196_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12147_ _09996_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12147_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12078_ _12077_/X _12446_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12078_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11029_ _11029_/A _11029_/B vssd1 vssd1 vccd1 vccd1 _12306_/D sky130_fd_sc_hd__nor2_1
XFILLER_77_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06570_ _06563_/X _06567_/X _06573_/A vssd1 vssd1 vccd1 vccd1 _06576_/A sky130_fd_sc_hd__a21oi_1
XFILLER_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08240_ _13106_/Q _08164_/Y _08239_/Y _12809_/Q vssd1 vssd1 vccd1 vccd1 _08240_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08171_ _13143_/Q _10482_/A _13127_/Q _10439_/A vssd1 vssd1 vccd1 vccd1 _08171_/X
+ sky130_fd_sc_hd__o22a_1
X_07122_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07122_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07053_ _07069_/A vssd1 vssd1 vccd1 vccd1 _07053_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07955_ _07961_/A vssd1 vssd1 vccd1 vccd1 _07955_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06906_ _06658_/A _06896_/X _06904_/X _06769_/A _06905_/Y vssd1 vssd1 vccd1 vccd1
+ _06907_/A sky130_fd_sc_hd__a32o_1
X_07886_ _12838_/Q vssd1 vssd1 vccd1 vccd1 _07886_/Y sky130_fd_sc_hd__inv_2
X_09625_ _09625_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09625_/Y sky130_fd_sc_hd__nand2_1
X_06837_ _06863_/A vssd1 vssd1 vccd1 vccd1 _06837_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09556_ _09524_/Y _09528_/A _09538_/A vssd1 vssd1 vccd1 vccd1 _09556_/Y sky130_fd_sc_hd__o21ai_2
X_06768_ _13201_/Q vssd1 vssd1 vccd1 vccd1 _06768_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08507_ _08518_/A vssd1 vssd1 vccd1 vccd1 _08507_/X sky130_fd_sc_hd__clkbuf_1
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06699_ _11987_/X _11990_/X _06698_/X vssd1 vssd1 vccd1 vccd1 _06699_/X sky130_fd_sc_hd__o21a_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09487_ _09487_/A vssd1 vssd1 vccd1 vccd1 _09490_/A sky130_fd_sc_hd__inv_2
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08438_ _08503_/A vssd1 vssd1 vccd1 vccd1 _08438_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_200_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08369_ _12799_/Q _08358_/X _07990_/X _08360_/X vssd1 vssd1 vccd1 vccd1 _12799_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10400_ _12924_/Q _10399_/Y _07809_/Y _10399_/A _10372_/X vssd1 vssd1 vccd1 vccd1
+ _10400_/X sky130_fd_sc_hd__o221a_1
X_11380_ _10590_/X _12404_/D _11404_/S vssd1 vssd1 vccd1 vccd1 _11380_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10331_ _10331_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _10333_/B sky130_fd_sc_hd__or2_4
XFILLER_139_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10262_ _13020_/Q _10228_/X _13053_/Q _10229_/X vssd1 vssd1 vccd1 vccd1 _10262_/X
+ sky130_fd_sc_hd__a22o_1
X_13050_ _12165_/X _13050_/D _07381_/X vssd1 vssd1 vccd1 vccd1 _13050_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12001_ _11063_/X _11062_/Y _12200_/S vssd1 vssd1 vccd1 vccd1 _12001_/X sky130_fd_sc_hd__mux2_1
X_10193_ _07881_/Y _10045_/A _08447_/Y _10113_/X vssd1 vssd1 vccd1 vccd1 _10193_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_160_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12903_ _12166_/X _12903_/D _07941_/X vssd1 vssd1 vccd1 vccd1 _12903_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12834_ _12169_/X _12834_/D _08282_/X vssd1 vssd1 vccd1 vccd1 _12834_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12765_/CLK _12765_/D _08509_/X vssd1 vssd1 vccd1 vccd1 _12765_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11716_ _11715_/X _10645_/Y _11774_/S vssd1 vssd1 vccd1 vccd1 _12422_/D sky130_fd_sc_hd__mux2_1
XPHY_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12696_ _12719_/CLK _12696_/D _08712_/X vssd1 vssd1 vccd1 vccd1 _12696_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _10517_/X _12932_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11647_/X sky130_fd_sc_hd__mux2_1
XPHY_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 io_in[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
XFILLER_30_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput24 io_in[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_1
Xinput35 io_in[6] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_1
XPHY_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput46 la_data_in[106] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_1
X_11578_ _12835_/Q _10793_/A _11578_/S vssd1 vssd1 vccd1 vccd1 _11578_/X sky130_fd_sc_hd__mux2_1
Xinput57 la_data_in[116] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_1
Xinput68 la_data_in[126] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_1
XFILLER_171_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10529_ _10529_/A _10529_/B _10529_/C vssd1 vssd1 vccd1 vccd1 _10529_/Y sky130_fd_sc_hd__nor3_4
XFILLER_7_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput79 la_data_in[20] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__buf_1
XFILLER_182_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13248_ _13249_/CLK _13248_/D _06378_/X vssd1 vssd1 vccd1 vccd1 _13248_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_131_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13179_ _13183_/CLK _13179_/D _06956_/X vssd1 vssd1 vccd1 vccd1 _13179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater614 _11610_/S vssd1 vssd1 vccd1 vccd1 _11603_/S sky130_fd_sc_hd__buf_6
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater625 _11578_/S vssd1 vssd1 vccd1 vccd1 _11569_/S sky130_fd_sc_hd__buf_4
X_07740_ _08556_/D _07750_/B vssd1 vssd1 vccd1 vccd1 _07740_/Y sky130_fd_sc_hd__nor2_1
Xrepeater636 input355/X vssd1 vssd1 vccd1 vccd1 _09186_/A sky130_fd_sc_hd__buf_8
Xrepeater647 _07980_/A vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__buf_8
XFILLER_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07671_ _07661_/A _07650_/B _07669_/X _07658_/B _07670_/X vssd1 vssd1 vccd1 vccd1
+ _07689_/D sky130_fd_sc_hd__o41a_1
XFILLER_26_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09410_ _12453_/Q _09384_/Y _12451_/Q _09418_/A _09409_/X vssd1 vssd1 vccd1 vccd1
+ _09422_/A sky130_fd_sc_hd__a221o_1
XFILLER_77_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06622_ _06650_/A vssd1 vssd1 vccd1 vccd1 _06622_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09341_ _12458_/Q vssd1 vssd1 vccd1 vccd1 _09341_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06553_ _06507_/X _06533_/Y _06489_/X _06552_/Y vssd1 vssd1 vccd1 vccd1 _13224_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_80_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09272_ _12303_/Q _12302_/Q vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__or2_1
X_06484_ _12044_/X _12043_/X _12044_/X _12043_/X vssd1 vssd1 vccd1 vccd1 _06484_/X
+ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_115_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 _12713_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08223_ _13104_/Q _10467_/B _13074_/Q vssd1 vssd1 vccd1 vccd1 _08238_/A sky130_fd_sc_hd__o21ai_1
XFILLER_20_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08154_ _12829_/Q vssd1 vssd1 vccd1 vccd1 _08154_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07105_ _07285_/A vssd1 vssd1 vccd1 vccd1 _07284_/A sky130_fd_sc_hd__inv_2
X_08085_ _08085_/A vssd1 vssd1 vccd1 vccd1 _08085_/X sky130_fd_sc_hd__clkbuf_1
X_07036_ _07735_/A vssd1 vssd1 vccd1 vccd1 _07069_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08987_ _12595_/Q vssd1 vssd1 vccd1 vccd1 _08995_/C sky130_fd_sc_hd__inv_2
XFILLER_130_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07938_ _12905_/Q _11494_/X _07946_/S vssd1 vssd1 vccd1 vccd1 _12905_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07869_ _13014_/Q vssd1 vssd1 vccd1 vccd1 _07869_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09608_ _09576_/Y _09592_/A _09589_/A vssd1 vssd1 vccd1 vccd1 _09608_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ _12336_/Q vssd1 vssd1 vccd1 vccd1 _10880_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09539_ _09524_/A _09524_/B _09538_/A _09524_/Y _09538_/Y vssd1 vssd1 vccd1 vccd1
+ _09555_/B sky130_fd_sc_hd__o32a_1
XFILLER_189_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12550_ _12550_/CLK _12550_/D _09068_/X vssd1 vssd1 vccd1 vccd1 _12550_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_185_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11501_ _10371_/Y input339/X _11501_/S vssd1 vssd1 vccd1 vccd1 _11501_/X sky130_fd_sc_hd__mux2_1
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12481_ _12485_/CLK _12481_/D vssd1 vssd1 vccd1 vccd1 _12481_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11432_ _12907_/Q _09243_/A _11443_/S vssd1 vssd1 vccd1 vccd1 _11432_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11363_ _12444_/Q _11362_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _11363_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13102_ _12167_/X _13102_/D _07230_/X vssd1 vssd1 vccd1 vccd1 _13102_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10314_ _13024_/Q _10049_/X _13057_/Q _10051_/X vssd1 vssd1 vccd1 vccd1 _10314_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11294_ vssd1 vssd1 vccd1 vccd1 _11294_/HI _11294_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13033_ _12164_/X _13033_/D _07433_/X vssd1 vssd1 vccd1 vccd1 _13033_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10245_ _10312_/A _11416_/X vssd1 vssd1 vccd1 vccd1 _10245_/Y sky130_fd_sc_hd__nor2b_4
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10176_ _13015_/Q _10049_/X _13048_/Q _10051_/X _10174_/X vssd1 vssd1 vccd1 vccd1
+ _10176_/X sky130_fd_sc_hd__a221o_1
XFILLER_78_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12817_ _12169_/X _12817_/D _08322_/X vssd1 vssd1 vccd1 vccd1 _12817_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12748_ _12749_/CLK _12748_/D _08581_/X vssd1 vssd1 vccd1 vccd1 _12748_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_187_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ _12679_/CLK _12679_/D _08762_/X vssd1 vssd1 vccd1 vccd1 _12679_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08910_ _08912_/A vssd1 vssd1 vccd1 vccd1 _08910_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_170_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09890_ _12655_/Q vssd1 vssd1 vccd1 vccd1 _09890_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08841_ _07746_/X _06278_/Y _08837_/X _12652_/Q vssd1 vssd1 vccd1 vccd1 _12652_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08772_ _08839_/A vssd1 vssd1 vccd1 vccd1 _08789_/A sky130_fd_sc_hd__clkbuf_2
X_07723_ _12948_/Q _07717_/X _07678_/A _07693_/X _07714_/X vssd1 vssd1 vccd1 vccd1
+ _12948_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07654_ _07654_/A _07654_/B _07690_/A vssd1 vssd1 vccd1 vccd1 _07676_/A sky130_fd_sc_hd__or3b_1
XFILLER_65_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06605_ _06605_/A vssd1 vssd1 vccd1 vccd1 _13219_/D sky130_fd_sc_hd__inv_2
XFILLER_41_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07585_ _12978_/Q _07574_/A _07568_/A _07575_/A _07583_/X vssd1 vssd1 vccd1 vccd1
+ _12978_/D sky130_fd_sc_hd__o221a_1
XFILLER_179_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09324_ _12365_/Q vssd1 vssd1 vccd1 vccd1 _09328_/A sky130_fd_sc_hd__inv_2
XFILLER_178_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06536_ _06982_/A vssd1 vssd1 vccd1 vccd1 _11083_/A sky130_fd_sc_hd__inv_2
XFILLER_179_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09255_ _12454_/Q _09250_/X _09244_/B _09251_/X vssd1 vssd1 vccd1 vccd1 _12454_/D
+ sky130_fd_sc_hd__a22o_1
X_06467_ _12765_/Q _12764_/Q vssd1 vssd1 vccd1 vccd1 _06468_/A sky130_fd_sc_hd__and2_1
X_08206_ _13091_/Q vssd1 vssd1 vccd1 vccd1 _08206_/Y sky130_fd_sc_hd__inv_2
X_09186_ _09186_/A _09186_/B _09186_/C _10558_/A vssd1 vssd1 vccd1 vccd1 _10535_/A
+ sky130_fd_sc_hd__or4_4
X_06398_ _06382_/X _12212_/X _06396_/X _06397_/X vssd1 vssd1 vccd1 vccd1 _13243_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08137_ _12824_/Q vssd1 vssd1 vccd1 vccd1 _10460_/A sky130_fd_sc_hd__inv_2
XFILLER_146_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08068_ _08083_/A vssd1 vssd1 vccd1 vccd1 _08068_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07019_ _07019_/A vssd1 vssd1 vccd1 vccd1 _11058_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10030_ _10027_/Y _10028_/X _10029_/Y _10134_/A vssd1 vssd1 vccd1 vccd1 _10041_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_103_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput203 la_oenb[17] vssd1 vssd1 vccd1 vccd1 input203/X sky130_fd_sc_hd__buf_1
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput214 la_oenb[27] vssd1 vssd1 vccd1 vccd1 input214/X sky130_fd_sc_hd__buf_1
Xinput225 la_oenb[37] vssd1 vssd1 vccd1 vccd1 input225/X sky130_fd_sc_hd__buf_1
XFILLER_89_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput236 la_oenb[47] vssd1 vssd1 vccd1 vccd1 input236/X sky130_fd_sc_hd__buf_1
XFILLER_88_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput247 la_oenb[57] vssd1 vssd1 vccd1 vccd1 input247/X sky130_fd_sc_hd__buf_1
Xinput258 la_oenb[67] vssd1 vssd1 vccd1 vccd1 input258/X sky130_fd_sc_hd__buf_1
Xinput269 la_oenb[77] vssd1 vssd1 vccd1 vccd1 input269/X sky130_fd_sc_hd__buf_1
XFILLER_5_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11981_ _10226_/Y _12797_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11981_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10932_ _10918_/Y _10919_/Y _10947_/A _10926_/X vssd1 vssd1 vccd1 vccd1 _10933_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10863_ _10861_/Y _10862_/Y _12522_/Q _12334_/Q vssd1 vssd1 vccd1 vccd1 _10890_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12602_ _12976_/CLK _12602_/D vssd1 vssd1 vccd1 vccd1 _12602_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10794_ _10794_/A _10794_/B _10794_/C _10794_/D vssd1 vssd1 vccd1 vccd1 _10795_/D
+ sky130_fd_sc_hd__or4_4
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12533_ _12537_/CLK _12533_/D vssd1 vssd1 vccd1 vccd1 _12533_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12464_ _12464_/CLK _12464_/D vssd1 vssd1 vccd1 vccd1 _12464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11415_ _10259_/Y _12799_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11415_/X sky130_fd_sc_hd__mux2_1
X_12395_ _12415_/CLK _12395_/D vssd1 vssd1 vccd1 vccd1 _12395_/Q sky130_fd_sc_hd__dfxtp_1
X_11346_ input39/X vssd1 vssd1 vccd1 vccd1 _11346_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11277_ vssd1 vssd1 vccd1 vccd1 _11277_/HI _11277_/LO sky130_fd_sc_hd__conb_1
X_13016_ _12164_/X _13016_/D _07473_/X vssd1 vssd1 vccd1 vccd1 _13016_/Q sky130_fd_sc_hd__dfrtp_1
X_10228_ _10276_/A vssd1 vssd1 vccd1 vccd1 _10228_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10159_ _10157_/Y _10000_/A _10158_/Y _10137_/X vssd1 vssd1 vccd1 vccd1 _10159_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07370_ _11431_/X _07368_/X _13055_/Q _07369_/X vssd1 vssd1 vccd1 vccd1 _13055_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06321_ _06105_/Y _06106_/Y _06108_/B _06320_/Y vssd1 vssd1 vccd1 vccd1 _06321_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_200_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06252_ _13273_/Q vssd1 vssd1 vccd1 vccd1 _06252_/Y sky130_fd_sc_hd__inv_2
X_09040_ _09071_/A _09267_/C _11967_/X _09433_/A vssd1 vssd1 vccd1 vccd1 _09043_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06183_ _06172_/A _06142_/Y _06136_/Y vssd1 vssd1 vccd1 vccd1 _06183_/X sky130_fd_sc_hd__o21a_1
XFILLER_190_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09942_ _09937_/Y _09922_/X _12045_/S _09938_/X _09941_/X vssd1 vssd1 vccd1 vccd1
+ _09942_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_132_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09873_ _13237_/Q vssd1 vssd1 vccd1 vccd1 _09873_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08824_ _08814_/X _08817_/X _06327_/Y _12659_/Q _08811_/X vssd1 vssd1 vccd1 vccd1
+ _12659_/D sky130_fd_sc_hd__a32o_1
X_08755_ _08769_/A vssd1 vssd1 vccd1 vccd1 _08755_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _12958_/Q _07694_/X _12957_/Q _07705_/X _07703_/X vssd1 vssd1 vccd1 vccd1
+ _12958_/D sky130_fd_sc_hd__o221a_1
XPHY_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08686_ _08686_/A vssd1 vssd1 vccd1 vccd1 _08686_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_130_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13264_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07637_ _12955_/Q _07646_/D _07637_/C vssd1 vssd1 vccd1 vccd1 _07637_/Y sky130_fd_sc_hd__nor3_4
XPHY_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07568_ _07568_/A vssd1 vssd1 vccd1 vccd1 _07568_/X sky130_fd_sc_hd__buf_4
XFILLER_201_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09307_ _08877_/X _07737_/X _07732_/X _12553_/Q _07037_/X vssd1 vssd1 vccd1 vccd1
+ _12553_/D sky130_fd_sc_hd__a41o_1
X_06519_ _06527_/A _06527_/B vssd1 vssd1 vccd1 vccd1 _06520_/B sky130_fd_sc_hd__and2_1
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07499_ _07778_/A vssd1 vssd1 vccd1 vccd1 _07522_/B sky130_fd_sc_hd__buf_2
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09238_ _12462_/Q _09231_/X _07562_/X _09233_/X vssd1 vssd1 vccd1 vccd1 _12462_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09169_ _11624_/X _09163_/X _12499_/Q _09164_/X vssd1 vssd1 vccd1 vccd1 _12499_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11200_ vssd1 vssd1 vccd1 vccd1 _11200_/HI _11200_/LO sky130_fd_sc_hd__conb_1
X_12180_ _10016_/X _12973_/Q _12180_/S vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11131_ _10730_/X _11075_/A _13253_/Q _11083_/A _12089_/X vssd1 vssd1 vccd1 vccd1
+ _11131_/X sky130_fd_sc_hd__a221o_1
XFILLER_89_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11062_ _11062_/A vssd1 vssd1 vccd1 vccd1 _11062_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10013_ _08739_/Y _10134_/A _06005_/Y _09972_/A _09991_/A vssd1 vssd1 vccd1 vccd1
+ _10013_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11964_ _12943_/Q _12941_/Q _11964_/S vssd1 vssd1 vccd1 vccd1 _11964_/X sky130_fd_sc_hd__mux2_1
X_10915_ _10915_/A vssd1 vssd1 vccd1 vccd1 _10921_/C sky130_fd_sc_hd__inv_2
XFILLER_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11895_ _10778_/X _10780_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _11895_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10846_ _10846_/A vssd1 vssd1 vccd1 vccd1 _10846_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10777_ _10763_/X _10768_/X _06379_/X _10769_/X _10770_/X vssd1 vssd1 vccd1 vccd1
+ _10777_/X sky130_fd_sc_hd__a221o_1
XFILLER_185_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12516_ _12849_/CLK _12516_/D vssd1 vssd1 vccd1 vccd1 _12516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12447_ _12492_/CLK _12447_/D vssd1 vssd1 vccd1 vccd1 _12447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput507 _11219_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput518 _11220_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12378_ _12577_/CLK _12378_/D vssd1 vssd1 vccd1 vccd1 _12400_/D sky130_fd_sc_hd__dfxtp_2
Xoutput529 _11221_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_125_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11329_ vssd1 vssd1 vccd1 vccd1 _11329_/HI _11329_/LO sky130_fd_sc_hd__conb_1
XFILLER_125_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06870_ _13189_/Q vssd1 vssd1 vccd1 vccd1 _06870_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08540_ _11962_/X _08562_/B vssd1 vssd1 vccd1 vccd1 _08541_/C sky130_fd_sc_hd__or2_1
XFILLER_82_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08471_ _13050_/Q vssd1 vssd1 vccd1 vccd1 _08471_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07422_ _07428_/A vssd1 vssd1 vccd1 vccd1 _07422_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07353_ _07368_/A vssd1 vssd1 vccd1 vccd1 _07353_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06304_ _06091_/B _06179_/Y _06090_/A _06179_/A vssd1 vssd1 vccd1 vccd1 _06305_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_149_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07284_ _07284_/A vssd1 vssd1 vccd1 vccd1 _11514_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_176_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09023_ _09023_/A input3/X vssd1 vssd1 vccd1 vccd1 _12575_/D sky130_fd_sc_hd__and2_1
X_06235_ _06245_/A vssd1 vssd1 vccd1 vccd1 _06235_/X sky130_fd_sc_hd__clkbuf_1
X_06166_ _07947_/A vssd1 vssd1 vccd1 vccd1 _08854_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06097_ _12726_/Q _12694_/Q _12726_/Q _12694_/Q vssd1 vssd1 vccd1 vccd1 _06098_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_160_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09925_ _12665_/Q vssd1 vssd1 vccd1 vccd1 _09925_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09856_ _06466_/Y _09844_/X _06462_/Y _09845_/X vssd1 vssd1 vccd1 vccd1 _09857_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_59_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08807_ _08807_/A vssd1 vssd1 vccd1 vccd1 _08807_/X sky130_fd_sc_hd__clkbuf_1
X_09787_ _06603_/Y _06607_/Y _09686_/A _09777_/Y vssd1 vssd1 vccd1 vccd1 _09787_/X
+ sky130_fd_sc_hd__o22a_1
X_06999_ _11852_/X vssd1 vssd1 vccd1 vccd1 _06999_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _08747_/A vssd1 vssd1 vccd1 vccd1 _08738_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _08669_/A vssd1 vssd1 vccd1 vccd1 _08669_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10700_ _06400_/X _10691_/A _10691_/B _10699_/X _10701_/A vssd1 vssd1 vccd1 vccd1
+ _10700_/X sky130_fd_sc_hd__a32o_1
XPHY_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11680_ _11679_/X _11380_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12382_/D sky130_fd_sc_hd__mux2_1
XPHY_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10631_ _10653_/B vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_14_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10562_ _10562_/A _10562_/B vssd1 vssd1 vccd1 vccd1 _10570_/A sky130_fd_sc_hd__nor2_4
XFILLER_167_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12301_ _12576_/CLK _12301_/D vssd1 vssd1 vccd1 vccd1 _12301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13281_ _13283_/CLK _13281_/D _06206_/X vssd1 vssd1 vccd1 vccd1 _13281_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10493_ _12498_/Q _09137_/B _09138_/B vssd1 vssd1 vccd1 vccd1 _10493_/X sky130_fd_sc_hd__a21bo_1
XFILLER_5_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12232_ _12231_/X _12636_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12232_/X sky130_fd_sc_hd__mux2_2
XFILLER_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _11146_/Y _10740_/X _12193_/S vssd1 vssd1 vccd1 vccd1 _12163_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11114_ _10686_/X _10737_/X _06410_/X _10738_/X _10739_/X vssd1 vssd1 vccd1 vccd1
+ _11114_/X sky130_fd_sc_hd__a221o_1
XFILLER_122_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12094_ _12448_/Q _12093_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12094_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11045_ _11045_/A vssd1 vssd1 vccd1 vccd1 _11045_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12996_ _12999_/CLK _12996_/D vssd1 vssd1 vccd1 vccd1 _12996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11947_ _09768_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11947_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11878_ _10313_/X _12819_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11878_/X sky130_fd_sc_hd__mux2_2
XFILLER_177_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10829_ _10828_/A _10828_/B _10827_/A _10827_/Y _10828_/Y vssd1 vssd1 vccd1 vccd1
+ _12328_/D sky130_fd_sc_hd__o32a_1
XFILLER_186_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06020_ _06272_/A vssd1 vssd1 vccd1 vccd1 _06314_/A sky130_fd_sc_hd__inv_2
XFILLER_142_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07971_ _11966_/X _10792_/C _09434_/B vssd1 vssd1 vccd1 vccd1 _08399_/B sky130_fd_sc_hd__or3_4
XFILLER_87_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09710_ _09708_/A _09708_/B _09709_/Y vssd1 vssd1 vccd1 vccd1 _09711_/B sky130_fd_sc_hd__a21o_1
X_06922_ _13183_/Q vssd1 vssd1 vccd1 vccd1 _09604_/B sky130_fd_sc_hd__inv_2
XFILLER_110_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09641_ _09641_/A vssd1 vssd1 vccd1 vccd1 _09641_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06853_ _06853_/A vssd1 vssd1 vccd1 vccd1 _06857_/A sky130_fd_sc_hd__inv_2
XFILLER_83_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09572_ _09572_/A _09572_/B vssd1 vssd1 vccd1 vccd1 _09574_/B sky130_fd_sc_hd__or2_2
X_06784_ _12034_/X vssd1 vssd1 vccd1 vccd1 _06785_/B sky130_fd_sc_hd__inv_2
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08523_ _08519_/X _12246_/X _08514_/X _12760_/Q vssd1 vssd1 vccd1 vccd1 _12760_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08454_ _13051_/Q vssd1 vssd1 vccd1 vccd1 _08454_/Y sky130_fd_sc_hd__inv_2
XPHY_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07405_ _08251_/A vssd1 vssd1 vccd1 vccd1 _08250_/A sky130_fd_sc_hd__inv_2
XFILLER_196_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08385_ _08385_/A vssd1 vssd1 vccd1 vccd1 _08385_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07336_ _11444_/X _07321_/X _13068_/Q _07324_/X vssd1 vssd1 vccd1 vccd1 _13068_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07267_ _11553_/X _07263_/X _13088_/Q _07264_/X vssd1 vssd1 vccd1 vccd1 _13088_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09006_ _09008_/A _09008_/B _11646_/X vssd1 vssd1 vccd1 vccd1 _12590_/D sky130_fd_sc_hd__and3_1
XFILLER_136_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06218_ _06046_/B _06210_/X _06046_/B _06210_/X vssd1 vssd1 vccd1 vccd1 _06218_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_117_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07198_ _08271_/A _10035_/A _09296_/A vssd1 vssd1 vccd1 vccd1 _11550_/S sky130_fd_sc_hd__nor3_4
XFILLER_3_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06149_ _12744_/Q _12712_/Q _06148_/X vssd1 vssd1 vccd1 vccd1 _06149_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09908_ _09906_/Y _09897_/X _06327_/A _09892_/X _09907_/X vssd1 vssd1 vccd1 vccd1
+ _09908_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_104_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09839_ _09839_/A _09839_/B vssd1 vssd1 vccd1 vccd1 _09839_/X sky130_fd_sc_hd__or2_2
XFILLER_132_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12850_ _12852_/CLK _12850_/D _08092_/X vssd1 vssd1 vccd1 vccd1 _12850_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _12065_/X _11800_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11801_/X sky130_fd_sc_hd__mux2_1
XPHY_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_12781_ _12852_/CLK _12781_/D _08416_/X vssd1 vssd1 vccd1 vccd1 _12781_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _09180_/D _11731_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11732_/X sky130_fd_sc_hd__mux2_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11383_/X _09185_/D _11675_/S vssd1 vssd1 vccd1 vccd1 _11663_/X sky130_fd_sc_hd__mux2_1
XPHY_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10614_ _11888_/S vssd1 vssd1 vccd1 vccd1 _10615_/B sky130_fd_sc_hd__inv_2
XPHY_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11594_ _10447_/Y _10528_/B _11603_/S vssd1 vssd1 vccd1 vccd1 _11594_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10545_ _12367_/Q _10541_/Y _09331_/B vssd1 vssd1 vccd1 vccd1 _10545_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_194_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13264_ _13264_/CLK _13264_/D _06302_/X vssd1 vssd1 vccd1 vccd1 _13264_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10476_ _10475_/A _10475_/B _10459_/X _10477_/B vssd1 vssd1 vccd1 vccd1 _10476_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12215_ _06323_/Y _13153_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12215_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13195_ _13196_/CLK _13195_/D _06828_/X vssd1 vssd1 vccd1 vccd1 _13195_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12146_ _09995_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12146_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12077_ _12446_/Q _12076_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12077_/X sky130_fd_sc_hd__mux2_1
X_11028_ _09150_/A _12305_/Q _09152_/A vssd1 vssd1 vccd1 vccd1 _11029_/B sky130_fd_sc_hd__o21a_1
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12979_ _12984_/CLK _12979_/D vssd1 vssd1 vccd1 vccd1 _12979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08170_ _10455_/B vssd1 vssd1 vccd1 vccd1 _10449_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07121_ _11544_/X _07113_/X _13143_/Q _07116_/X vssd1 vssd1 vccd1 vccd1 _13143_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07052_ _07063_/A vssd1 vssd1 vccd1 vccd1 _07052_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07954_ _12899_/Q _11488_/X _07962_/S vssd1 vssd1 vccd1 vccd1 _12899_/D sky130_fd_sc_hd__mux2_1
X_06905_ _13186_/Q vssd1 vssd1 vccd1 vccd1 _06905_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07885_ _12837_/Q vssd1 vssd1 vccd1 vccd1 _07885_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09624_ _09625_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09624_/X sky130_fd_sc_hd__or2_1
X_06836_ _06829_/X _06830_/Y _06769_/X _06835_/X vssd1 vssd1 vccd1 vccd1 _13195_/D
+ sky130_fd_sc_hd__o22ai_1
X_09555_ _09555_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09574_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_37_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12369_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_06767_ _06806_/A vssd1 vssd1 vccd1 vccd1 _06767_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08506_ _08521_/A vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_197_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09486_ _09471_/X _09487_/A _09483_/Y _09485_/X vssd1 vssd1 vccd1 vccd1 _09486_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_180_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06698_ _11986_/X _06698_/B vssd1 vssd1 vccd1 vccd1 _06698_/X sky130_fd_sc_hd__or2_2
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08437_ _12773_/Q _08417_/A _07566_/X _08418_/A vssd1 vssd1 vccd1 vccd1 _12773_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08368_ _08370_/A vssd1 vssd1 vccd1 vccd1 _08368_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07319_ _12843_/Q _11433_/S vssd1 vssd1 vccd1 vccd1 _07384_/A sky130_fd_sc_hd__or2_2
XFILLER_178_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08299_ _08372_/A vssd1 vssd1 vccd1 vccd1 _08311_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10330_ _10328_/A _10328_/B _10329_/Y _10324_/A vssd1 vssd1 vccd1 vccd1 _10330_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_192_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ _13093_/Q _10228_/X _13125_/Q _10229_/X vssd1 vssd1 vccd1 vccd1 _10261_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12000_ _11078_/X _11069_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12000_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10192_ _08199_/Y _10151_/X _10191_/X vssd1 vssd1 vccd1 vccd1 _10192_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12902_ _12166_/X _12902_/D _07943_/X vssd1 vssd1 vccd1 vccd1 _12902_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12833_ _12169_/X _12833_/D _08285_/X vssd1 vssd1 vccd1 vccd1 _12833_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12764_ _12769_/CLK _12764_/D _08511_/X vssd1 vssd1 vccd1 vccd1 _12764_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _10645_/Y _10646_/Y _11818_/S vssd1 vssd1 vccd1 vccd1 _11715_/X sky130_fd_sc_hd__mux2_1
XPHY_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12695_ _12695_/CLK _12695_/D _08714_/X vssd1 vssd1 vccd1 vccd1 _12695_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_159_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11646_ _10516_/X _12931_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11646_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 io_in[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_1
XFILLER_35_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput25 io_in[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_1
XPHY_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput36 io_in[7] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_1
XPHY_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11577_ _12834_/Q _10793_/B _11578_/S vssd1 vssd1 vccd1 vccd1 _11577_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput47 la_data_in[107] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_1
Xinput58 la_data_in[117] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_1
X_10528_ _10528_/A _10528_/B _10528_/C _09243_/A vssd1 vssd1 vccd1 vccd1 _10529_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_7_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput69 la_data_in[127] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_1
XFILLER_183_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13247_ _13249_/CLK _13247_/D _06381_/X vssd1 vssd1 vccd1 vccd1 _13247_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_171_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10459_ _10459_/A vssd1 vssd1 vccd1 vccd1 _10459_/X sky130_fd_sc_hd__buf_2
XFILLER_124_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13178_ _13183_/CLK _13178_/D _06973_/X vssd1 vssd1 vccd1 vccd1 _13178_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12129_ _12128_/X _12437_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12129_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater615 _08271_/Y vssd1 vssd1 vccd1 vccd1 _11610_/S sky130_fd_sc_hd__buf_6
Xrepeater626 _11550_/S vssd1 vssd1 vccd1 vccd1 _11578_/S sky130_fd_sc_hd__buf_4
Xrepeater637 input354/X vssd1 vssd1 vccd1 vccd1 _09186_/B sky130_fd_sc_hd__buf_8
XFILLER_65_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater648 input333/X vssd1 vssd1 vccd1 vccd1 _10528_/C sky130_fd_sc_hd__buf_8
X_07670_ _07678_/A _12946_/Q _07670_/C _12948_/Q vssd1 vssd1 vccd1 vccd1 _07670_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_93_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06621_ _06507_/X _06607_/Y _06608_/X _06620_/Y vssd1 vssd1 vccd1 vccd1 _13218_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_19_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09340_ _09335_/Y _12397_/Q _09336_/Y _12404_/Q _09339_/X vssd1 vssd1 vccd1 vccd1
+ _09340_/X sky130_fd_sc_hd__a221o_1
XFILLER_179_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06552_ _06552_/A _06552_/B vssd1 vssd1 vccd1 vccd1 _06552_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09271_ _09271_/A _12301_/Q _09271_/C vssd1 vssd1 vccd1 vccd1 _09271_/X sky130_fd_sc_hd__and3_1
XFILLER_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06483_ _13230_/Q vssd1 vssd1 vccd1 vccd1 _06483_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08222_ _08222_/A _08222_/B _08219_/X _08221_/X vssd1 vssd1 vccd1 vccd1 _08247_/B
+ sky130_fd_sc_hd__or4bb_4
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08153_ _13141_/Q _10477_/A _08129_/Y _12813_/Q vssd1 vssd1 vccd1 vccd1 _08153_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_155_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12751_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07104_ _08271_/A _10090_/A _09296_/A vssd1 vssd1 vccd1 vccd1 _07285_/A sky130_fd_sc_hd__or3_4
XFILLER_147_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08084_ _12854_/Q _08082_/X _07997_/X _08083_/X vssd1 vssd1 vccd1 vccd1 _12854_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07035_ _12613_/Q vssd1 vssd1 vccd1 vccd1 _07735_/A sky130_fd_sc_hd__buf_2
XFILLER_103_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08986_ _09283_/A _08986_/B vssd1 vssd1 vccd1 vccd1 _12601_/D sky130_fd_sc_hd__nor2_1
XFILLER_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07937_ _07945_/A vssd1 vssd1 vccd1 vccd1 _07937_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07868_ _12917_/Q vssd1 vssd1 vccd1 vccd1 _07868_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06819_ _06817_/X _06818_/X _06817_/X _06818_/X vssd1 vssd1 vccd1 vccd1 _06819_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_09607_ _09607_/A _09607_/B vssd1 vssd1 vccd1 vccd1 _09632_/A sky130_fd_sc_hd__or2_1
XFILLER_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07799_ _13012_/Q vssd1 vssd1 vccd1 vccd1 _07799_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09538_ _09538_/A vssd1 vssd1 vccd1 vccd1 _09538_/Y sky130_fd_sc_hd__inv_2
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09469_ _09469_/A vssd1 vssd1 vccd1 vccd1 _11958_/S sky130_fd_sc_hd__inv_16
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11500_ _10366_/X input338/X _11501_/S vssd1 vssd1 vccd1 vccd1 _11500_/X sky130_fd_sc_hd__mux2_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12480_ _12480_/CLK _12480_/D vssd1 vssd1 vccd1 vccd1 _12480_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11431_ _12906_/Q _10528_/C _11433_/S vssd1 vssd1 vccd1 vccd1 _11431_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11362_ _12444_/Q _10660_/Y _12091_/S vssd1 vssd1 vccd1 vccd1 _11362_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13101_ _12167_/X _13101_/D _07232_/X vssd1 vssd1 vccd1 vccd1 _13101_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10313_ _13097_/Q _10049_/X _13129_/Q _10051_/X vssd1 vssd1 vccd1 vccd1 _10313_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11293_ vssd1 vssd1 vccd1 vccd1 _11293_/HI _11293_/LO sky130_fd_sc_hd__conb_1
X_13032_ _12164_/X _13032_/D _07435_/X vssd1 vssd1 vccd1 vccd1 _13032_/Q sky130_fd_sc_hd__dfrtp_1
X_10244_ _10244_/A vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__buf_6
XFILLER_106_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10175_ _13088_/Q _10049_/X _13120_/Q _10051_/X _10174_/X vssd1 vssd1 vccd1 vccd1
+ _10175_/X sky130_fd_sc_hd__a221o_1
XFILLER_191_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12816_ _12169_/X _12816_/D _08325_/X vssd1 vssd1 vccd1 vccd1 _12816_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12747_ _12747_/CLK _12747_/D _08583_/X vssd1 vssd1 vccd1 vccd1 _12747_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_163_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _12679_/CLK _12678_/D _08766_/X vssd1 vssd1 vccd1 vccd1 _12678_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_187_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11629_ _10499_/X _12928_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11629_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08840_ _08851_/A vssd1 vssd1 vccd1 vccd1 _08840_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08771_ _08770_/Y _08760_/X _06228_/X _08764_/X vssd1 vssd1 vccd1 vccd1 _12677_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_100_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07722_ _12949_/Q _07717_/X _12948_/Q _07693_/X _07714_/X vssd1 vssd1 vccd1 vccd1
+ _12949_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07653_ _07649_/Y _12950_/Q _07651_/B _08980_/A _07652_/X vssd1 vssd1 vccd1 vccd1
+ _07690_/A sky130_fd_sc_hd__o311a_1
XFILLER_93_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06604_ _06526_/X _06598_/B _06602_/Y _06556_/X _06603_/Y vssd1 vssd1 vccd1 vccd1
+ _06605_/A sky130_fd_sc_hd__o32a_1
XFILLER_129_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07584_ _12979_/Q _07574_/A _09226_/B _07575_/A _07583_/X vssd1 vssd1 vccd1 vccd1
+ _12979_/D sky130_fd_sc_hd__o221a_1
X_09323_ _12366_/Q vssd1 vssd1 vccd1 vccd1 _09329_/A sky130_fd_sc_hd__inv_2
XFILLER_179_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06535_ _06535_/A _12762_/Q vssd1 vssd1 vccd1 vccd1 _06982_/A sky130_fd_sc_hd__or2b_2
XFILLER_178_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09254_ _12455_/Q _09250_/X _09244_/A _09251_/X vssd1 vssd1 vccd1 vccd1 _12455_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06466_ _13232_/Q vssd1 vssd1 vccd1 vccd1 _06466_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08205_ _13103_/Q vssd1 vssd1 vccd1 vccd1 _08205_/Y sky130_fd_sc_hd__inv_2
X_09185_ _09185_/A _09185_/B _09185_/C _09185_/D vssd1 vssd1 vccd1 vccd1 _10558_/A
+ sky130_fd_sc_hd__or4_4
X_06397_ _13243_/Q vssd1 vssd1 vccd1 vccd1 _06397_/X sky130_fd_sc_hd__buf_2
XFILLER_105_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08136_ _12809_/Q vssd1 vssd1 vccd1 vccd1 _10418_/A sky130_fd_sc_hd__inv_2
XFILLER_105_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08067_ _08067_/A vssd1 vssd1 vccd1 vccd1 _08083_/A sky130_fd_sc_hd__inv_2
XFILLER_49_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07018_ _07024_/A vssd1 vssd1 vccd1 vccd1 _07018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput204 la_oenb[18] vssd1 vssd1 vccd1 vccd1 input204/X sky130_fd_sc_hd__buf_1
XFILLER_49_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput215 la_oenb[28] vssd1 vssd1 vccd1 vccd1 input215/X sky130_fd_sc_hd__buf_1
Xinput226 la_oenb[38] vssd1 vssd1 vccd1 vccd1 input226/X sky130_fd_sc_hd__buf_1
Xinput237 la_oenb[48] vssd1 vssd1 vccd1 vccd1 input237/X sky130_fd_sc_hd__buf_1
XFILLER_76_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13004_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput248 la_oenb[58] vssd1 vssd1 vccd1 vccd1 input248/X sky130_fd_sc_hd__buf_1
XFILLER_75_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput259 la_oenb[68] vssd1 vssd1 vccd1 vccd1 input259/X sky130_fd_sc_hd__buf_1
X_08969_ _08969_/A vssd1 vssd1 vccd1 vccd1 _08969_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11980_ _10206_/Y _12796_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10931_ _10930_/A _10930_/B _10930_/Y vssd1 vssd1 vccd1 vccd1 _10934_/A sky130_fd_sc_hd__a21oi_2
XFILLER_112_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ _12334_/Q vssd1 vssd1 vccd1 vccd1 _10862_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12977_/CLK _12601_/D vssd1 vssd1 vccd1 vccd1 _12601_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _10793_/A _10793_/B vssd1 vssd1 vccd1 vccd1 _10795_/C sky130_fd_sc_hd__or2_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12532_ _12537_/CLK _12532_/D vssd1 vssd1 vccd1 vccd1 _12532_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_200_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12463_ _12985_/CLK _12463_/D vssd1 vssd1 vccd1 vccd1 _12463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11414_ _11413_/X _12443_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _11414_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12394_ _12467_/CLK _12394_/D vssd1 vssd1 vccd1 vccd1 _12416_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11345_ _11345_/A vssd1 vssd1 vccd1 vccd1 _11345_/X sky130_fd_sc_hd__buf_1
XFILLER_153_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11276_ vssd1 vssd1 vccd1 vccd1 _11276_/HI _11276_/LO sky130_fd_sc_hd__conb_1
XFILLER_140_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13015_ _12164_/X _13015_/D _07479_/X vssd1 vssd1 vccd1 vccd1 _13015_/Q sky130_fd_sc_hd__dfrtp_2
X_10227_ _10227_/A _11981_/X vssd1 vssd1 vccd1 vccd1 _10227_/Y sky130_fd_sc_hd__nor2b_4
X_10158_ _12851_/Q vssd1 vssd1 vccd1 vccd1 _10158_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10089_ _10150_/A _11974_/X vssd1 vssd1 vccd1 vccd1 _10089_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_48_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06320_ _06320_/A vssd1 vssd1 vccd1 vccd1 _06320_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06251_ _06280_/A vssd1 vssd1 vccd1 vccd1 _06251_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06182_ _06182_/A _06182_/B _06209_/C vssd1 vssd1 vccd1 vccd1 _06182_/X sky130_fd_sc_hd__or3_2
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09941_ _09941_/A vssd1 vssd1 vccd1 vccd1 _09941_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09872_ _09492_/X _09870_/Y _09877_/A _09700_/A vssd1 vssd1 vccd1 vccd1 _09872_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_112_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08823_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08823_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08754_ _08753_/Y _08565_/X _06200_/X _08742_/X vssd1 vssd1 vccd1 vccd1 _12682_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _07705_/A vssd1 vssd1 vccd1 vccd1 _07705_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _08685_/A vssd1 vssd1 vccd1 vccd1 _08685_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _12957_/Q _12956_/Q _07665_/B _07664_/A vssd1 vssd1 vccd1 vccd1 _07637_/C
+ sky130_fd_sc_hd__or4_4
XPHY_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07567_ _07566_/X _07552_/A _12987_/Q _07553_/A _07556_/X vssd1 vssd1 vccd1 vccd1
+ _12987_/D sky130_fd_sc_hd__a221o_1
XFILLER_94_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09306_ _08877_/X _07737_/X _07732_/X _12617_/Q _08908_/X vssd1 vssd1 vccd1 vccd1
+ _12617_/D sky130_fd_sc_hd__a41o_1
X_06518_ _12042_/X _06497_/A _06495_/Y _06497_/Y vssd1 vssd1 vccd1 vccd1 _06527_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_194_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07498_ _09267_/C _12312_/Q vssd1 vssd1 vccd1 vccd1 _07778_/A sky130_fd_sc_hd__nand2_4
XFILLER_181_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09237_ _12463_/Q _09231_/X _07560_/X _09233_/X vssd1 vssd1 vccd1 vccd1 _12463_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06449_ _06356_/X _06860_/A _06427_/X _10711_/A _06448_/Y vssd1 vssd1 vccd1 vccd1
+ _06451_/A sky130_fd_sc_hd__o221a_2
XFILLER_182_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09168_ _11625_/X _09163_/X _12500_/Q _09164_/X vssd1 vssd1 vccd1 vccd1 _12500_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08119_ _08112_/Y _08113_/X _08114_/Y _10475_/A _08118_/X vssd1 vssd1 vccd1 vccd1
+ _08132_/B sky130_fd_sc_hd__a221o_1
XFILLER_181_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09099_ _09115_/A vssd1 vssd1 vccd1 vccd1 _09099_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11130_ _11041_/A _10788_/X _13244_/Q _11111_/X _11112_/X vssd1 vssd1 vccd1 vccd1
+ _11130_/X sky130_fd_sc_hd__a221o_1
XFILLER_79_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11061_ _11033_/X _11054_/X _06397_/X _11055_/X _11060_/X vssd1 vssd1 vccd1 vccd1
+ _11061_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10012_ _08745_/Y _10134_/A _06169_/Y _09972_/A _09991_/A vssd1 vssd1 vccd1 vccd1
+ _10012_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_95_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11963_ _06025_/B _06025_/A _11963_/S vssd1 vssd1 vccd1 vccd1 _11963_/X sky130_fd_sc_hd__mux2_2
XFILLER_44_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10914_ _12528_/Q _12340_/Q _10908_/X _10909_/X vssd1 vssd1 vccd1 vccd1 _10916_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11894_ _10777_/X _10771_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _11894_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10845_ _10837_/Y _10838_/Y _10836_/Y _10864_/A vssd1 vssd1 vccd1 vccd1 _10846_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10776_ _10755_/X _10759_/X _06371_/X _10760_/X _10761_/X vssd1 vssd1 vccd1 vccd1
+ _10776_/X sky130_fd_sc_hd__a221o_1
X_12515_ _12849_/CLK _12515_/D vssd1 vssd1 vccd1 vccd1 _12515_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_121_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12446_ _12492_/CLK _12446_/D vssd1 vssd1 vccd1 vccd1 _12446_/Q sky130_fd_sc_hd__dfxtp_1
X_12377_ _12577_/CLK _12377_/D vssd1 vssd1 vccd1 vccd1 _12399_/D sky130_fd_sc_hd__dfxtp_2
Xoutput508 _11256_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__clkbuf_2
Xoutput519 _11266_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ vssd1 vssd1 vccd1 vccd1 _11328_/HI _11328_/LO sky130_fd_sc_hd__conb_1
XFILLER_181_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11259_ vssd1 vssd1 vccd1 vccd1 _11259_/HI _11259_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08470_ _13060_/Q _10367_/B _13053_/Q _10346_/A vssd1 vssd1 vccd1 vccd1 _08473_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_91_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07421_ _11479_/X _07412_/X _13038_/Q _07415_/X vssd1 vssd1 vccd1 vccd1 _13038_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_196_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07352_ _07360_/A vssd1 vssd1 vccd1 vccd1 _07352_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_188_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06303_ _12608_/Q vssd1 vssd1 vccd1 vccd1 _06303_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_176_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07283_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07283_/X sky130_fd_sc_hd__clkbuf_1
X_09022_ _09023_/A _12575_/Q vssd1 vssd1 vccd1 vccd1 _12576_/D sky130_fd_sc_hd__and2_1
XFILLER_176_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06234_ _06231_/Y _06216_/X _06217_/X _06233_/X vssd1 vssd1 vccd1 vccd1 _13277_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_164_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06165_ _07590_/A vssd1 vssd1 vccd1 vccd1 _07947_/A sky130_fd_sc_hd__inv_2
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _12328_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06096_ _12728_/Q _12696_/Q _06095_/X vssd1 vssd1 vccd1 vccd1 _06096_/X sky130_fd_sc_hd__o21a_1
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09924_ _09921_/Y _09922_/X _06300_/A _09915_/X _09923_/X vssd1 vssd1 vccd1 vccd1
+ _09924_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_160_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09855_ _09492_/X _09853_/Y _09860_/A _09700_/A vssd1 vssd1 vccd1 vccd1 _09855_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08806_ _08798_/X _08801_/X _06291_/Y _12666_/Q _08567_/X vssd1 vssd1 vccd1 vccd1
+ _12666_/D sky130_fd_sc_hd__a32o_1
XFILLER_105_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09786_ _09701_/X _09784_/Y _09785_/X _09682_/X vssd1 vssd1 vccd1 vccd1 _09786_/X
+ sky130_fd_sc_hd__a31o_1
X_06998_ _13173_/Q vssd1 vssd1 vccd1 vccd1 _09524_/B sky130_fd_sc_hd__inv_2
XFILLER_86_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08737_ _11820_/X _08592_/A _12686_/Q _08593_/A vssd1 vssd1 vccd1 vccd1 _12686_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _11848_/X _08654_/X _12714_/Q _08655_/X vssd1 vssd1 vccd1 vccd1 _12714_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ _11612_/X _07610_/A _12967_/Q _07611_/A _07616_/X vssd1 vssd1 vccd1 vccd1
+ _12967_/D sky130_fd_sc_hd__o221a_1
XFILLER_14_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _11950_/X _08592_/X _12741_/Q _08593_/X vssd1 vssd1 vccd1 vccd1 _12741_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _12103_/S _10796_/D vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__or2_1
XPHY_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ _10561_/A vssd1 vssd1 vccd1 vccd1 _10562_/B sky130_fd_sc_hd__inv_2
XFILLER_194_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12300_ _12576_/CLK _12300_/D vssd1 vssd1 vccd1 vccd1 _12300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13280_ _13283_/CLK _13280_/D _06214_/X vssd1 vssd1 vccd1 vccd1 _13280_/Q sky130_fd_sc_hd__dfrtp_1
X_10492_ _12497_/Q _09136_/B _09137_/B vssd1 vssd1 vccd1 vccd1 _10492_/X sky130_fd_sc_hd__a21bo_1
XFILLER_108_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12231_ _06278_/Y _13161_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12231_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12162_ _11145_/Y _11144_/X _12193_/S vssd1 vssd1 vccd1 vccd1 _12162_/X sky130_fd_sc_hd__mux2_2
XFILLER_162_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11113_ _10696_/X _10788_/X _13241_/Q _11111_/X _11112_/X vssd1 vssd1 vccd1 vccd1
+ _11113_/X sky130_fd_sc_hd__a221o_1
XFILLER_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12093_ _12092_/X _12448_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12093_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11044_ _10693_/X _10746_/X _06407_/X _07008_/X _10747_/X vssd1 vssd1 vccd1 vccd1
+ _11044_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12995_ _12995_/CLK _12995_/D vssd1 vssd1 vccd1 vccd1 _12995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11946_ _09754_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11946_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11877_ _10308_/X _12818_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11877_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10828_ _10828_/A _10828_/B vssd1 vssd1 vccd1 vccd1 _10828_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ _10759_/A vssd1 vssd1 vccd1 vccd1 _10759_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_187_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12429_ _12474_/CLK _12429_/D vssd1 vssd1 vccd1 vccd1 _12429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07970_ _12549_/Q vssd1 vssd1 vccd1 vccd1 _10792_/C sky130_fd_sc_hd__inv_2
XFILLER_113_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06921_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06921_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06852_ _12025_/X _12021_/X _06846_/X _06847_/X _06851_/X vssd1 vssd1 vccd1 vccd1
+ _06853_/A sky130_fd_sc_hd__o32a_1
XFILLER_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09640_ _09640_/A _09640_/B vssd1 vssd1 vccd1 vccd1 _09641_/A sky130_fd_sc_hd__or2_1
XFILLER_132_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_109_wb_clk_i _12726_/CLK vssd1 vssd1 vccd1 vccd1 _12737_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09571_ _09471_/X _09567_/X _09568_/Y _09570_/X vssd1 vssd1 vccd1 vccd1 _09571_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_167_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06783_ _06783_/A _06783_/B vssd1 vssd1 vccd1 vccd1 _06783_/X sky130_fd_sc_hd__or2_1
XFILLER_67_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08522_ _08533_/A vssd1 vssd1 vccd1 vccd1 _08522_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ _13063_/Q vssd1 vssd1 vccd1 vccd1 _08453_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07404_ _08271_/A _10090_/A _09295_/A vssd1 vssd1 vccd1 vccd1 _08251_/A sky130_fd_sc_hd__or3_4
XPHY_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08384_ _12793_/Q _08374_/X _07293_/X _08375_/X vssd1 vssd1 vccd1 vccd1 _12793_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07335_ _07345_/A vssd1 vssd1 vccd1 vccd1 _07335_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07266_ _07266_/A vssd1 vssd1 vccd1 vccd1 _07266_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09005_ _09008_/A _09008_/B _11647_/X vssd1 vssd1 vccd1 vccd1 _12591_/D sky130_fd_sc_hd__and3_1
XFILLER_191_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06217_ _06217_/A vssd1 vssd1 vccd1 vccd1 _06217_/X sky130_fd_sc_hd__clkbuf_2
X_07197_ _09976_/B vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06148_ _12744_/Q _12712_/Q _12743_/Q _12711_/Q vssd1 vssd1 vccd1 vccd1 _06148_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06079_ _12732_/Q _12700_/Q _06078_/X vssd1 vssd1 vccd1 vccd1 _06079_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_104_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09907_ _12882_/Q _09910_/B vssd1 vssd1 vccd1 vccd1 _09907_/X sky130_fd_sc_hd__or2_1
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09838_ _13231_/Q _09837_/A _09836_/Y _09837_/Y vssd1 vssd1 vccd1 vccd1 _09839_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09769_ _09769_/A _09769_/B vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _10528_/B _11799_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11800_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12780_ _12852_/CLK _12780_/D _08420_/X vssd1 vssd1 vccd1 vccd1 _12780_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11414_/X _12487_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11731_/X sky130_fd_sc_hd__mux2_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11661_/X _11384_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12373_/D sky130_fd_sc_hd__mux2_1
XPHY_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ _11406_/X vssd1 vssd1 vccd1 vccd1 _10625_/A sky130_fd_sc_hd__inv_2
XPHY_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11593_ _10443_/X _09243_/A _11603_/S vssd1 vssd1 vccd1 vccd1 _11593_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10544_ _11359_/X _10554_/B vssd1 vssd1 vccd1 vccd1 _10544_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13263_ _13264_/CLK _13263_/D _06308_/X vssd1 vssd1 vccd1 vccd1 _13263_/Q sky130_fd_sc_hd__dfrtp_1
X_10475_ _10475_/A _10475_/B vssd1 vssd1 vccd1 vccd1 _10477_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12214_ _12213_/X _12627_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12214_/X sky130_fd_sc_hd__mux2_2
X_13194_ _13237_/CLK _13194_/D _06837_/X vssd1 vssd1 vccd1 vccd1 _13194_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12145_ _09994_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12145_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_7_wb_clk_i _12328_/CLK vssd1 vssd1 vccd1 vccd1 _12868_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12076_ _12075_/X _12446_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12076_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11027_ _08191_/X _08275_/Y _13079_/Q vssd1 vssd1 vccd1 vccd1 _12554_/D sky130_fd_sc_hd__o21a_1
XFILLER_38_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12978_ _12978_/CLK _12978_/D vssd1 vssd1 vccd1 vccd1 _12978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11929_ _09496_/Y _12790_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11929_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07120_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07120_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07051_ _07037_/X _07040_/X _06291_/Y _13159_/Q _07042_/X vssd1 vssd1 vccd1 vccd1
+ _13159_/D sky130_fd_sc_hd__a32o_1
XFILLER_103_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07953_ _07961_/A vssd1 vssd1 vccd1 vccd1 _07953_/X sky130_fd_sc_hd__clkbuf_1
X_06904_ _12024_/X _12020_/X _06898_/X _06899_/X _06903_/X vssd1 vssd1 vccd1 vccd1
+ _06904_/X sky130_fd_sc_hd__o32a_2
XFILLER_29_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07884_ _08271_/A _09969_/B _09295_/A vssd1 vssd1 vccd1 vccd1 _11487_/S sky130_fd_sc_hd__nor3_4
XFILLER_68_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ _09630_/A _09623_/B vssd1 vssd1 vccd1 vccd1 _09625_/B sky130_fd_sc_hd__or2_1
X_06835_ _06831_/X _06832_/X _06821_/X _06813_/X _06834_/X vssd1 vssd1 vccd1 vccd1
+ _06835_/X sky130_fd_sc_hd__o221a_1
XFILLER_55_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06766_ _06766_/A vssd1 vssd1 vccd1 vccd1 _06806_/A sky130_fd_sc_hd__clkbuf_2
X_09554_ _09566_/A _09554_/B vssd1 vssd1 vccd1 vccd1 _09572_/A sky130_fd_sc_hd__or2_1
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08505_ _08504_/X _12260_/X _08499_/X _12767_/Q vssd1 vssd1 vccd1 vccd1 _12767_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09485_ _09484_/Y _07735_/A _12862_/Q _07729_/X vssd1 vssd1 vccd1 vccd1 _09485_/X
+ sky130_fd_sc_hd__a22o_1
X_06697_ _13254_/Q _10687_/A _12755_/Q _06427_/A _11034_/A vssd1 vssd1 vccd1 vccd1
+ _06698_/B sky130_fd_sc_hd__a32o_1
XFILLER_197_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08436_ _08503_/A vssd1 vssd1 vccd1 vccd1 _08436_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_77_wb_clk_i _13219_/CLK vssd1 vssd1 vccd1 vccd1 _13196_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08367_ _12800_/Q _08358_/X _07986_/X _08360_/X vssd1 vssd1 vccd1 vccd1 _12800_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07318_ _07409_/A _09978_/B _09295_/A vssd1 vssd1 vccd1 vccd1 _11422_/S sky130_fd_sc_hd__nor3_4
XFILLER_176_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08298_ _08657_/A vssd1 vssd1 vccd1 vccd1 _08372_/A sky130_fd_sc_hd__buf_6
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07249_ _07249_/A vssd1 vssd1 vccd1 vccd1 _07249_/X sky130_fd_sc_hd__buf_2
XFILLER_109_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10260_ _10312_/A _11415_/X vssd1 vssd1 vccd1 vccd1 _10260_/Y sky130_fd_sc_hd__nor2b_4
XFILLER_124_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10191_ _08269_/Y _10045_/A _08116_/Y _10113_/X vssd1 vssd1 vccd1 vccd1 _10191_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12901_ _12166_/X _12901_/D _07945_/X vssd1 vssd1 vccd1 vccd1 _12901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12832_ _12169_/X _12832_/D _08287_/X vssd1 vssd1 vccd1 vccd1 _12832_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12763_ _12773_/CLK _12763_/D _08513_/X vssd1 vssd1 vccd1 vccd1 _12763_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11714_ _11713_/X _10641_/Y _11774_/S vssd1 vssd1 vccd1 vccd1 _12421_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12695_/CLK _12694_/D _08719_/X vssd1 vssd1 vccd1 vccd1 _12694_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _10515_/X _12930_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11645_/X sky130_fd_sc_hd__mux2_1
XPHY_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 io_in[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_1
Xinput26 io_in[32] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
XFILLER_35_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11576_ _12833_/Q _10794_/A _11578_/S vssd1 vssd1 vccd1 vccd1 _11576_/X sky130_fd_sc_hd__mux2_1
Xinput37 io_in[8] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_1
XPHY_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput48 la_data_in[108] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_1
XFILLER_128_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput59 la_data_in[118] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_1
XFILLER_182_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10527_ _10527_/A _10527_/B _10527_/C _10527_/D vssd1 vssd1 vccd1 vccd1 _11704_/S
+ sky130_fd_sc_hd__or4_4
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13246_ _13249_/CLK _13246_/D _06385_/X vssd1 vssd1 vccd1 vccd1 _13246_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_108_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10458_ _10458_/A _10463_/C _10458_/C vssd1 vssd1 vccd1 vccd1 _10458_/Y sky130_fd_sc_hd__nor3_1
XFILLER_6_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10389_ _10388_/A _10388_/B _10372_/X _10390_/B vssd1 vssd1 vccd1 vccd1 _10389_/X
+ sky130_fd_sc_hd__o211a_1
X_13177_ _13177_/CLK _13177_/D _06976_/X vssd1 vssd1 vccd1 vccd1 _13177_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12128_ _12437_/Q _12127_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12128_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12059_ _12058_/X _12439_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12059_/X sky130_fd_sc_hd__mux2_1
Xrepeater616 _11501_/S vssd1 vssd1 vccd1 vccd1 _11513_/S sky130_fd_sc_hd__buf_6
XFILLER_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater627 _11550_/S vssd1 vssd1 vccd1 vccd1 _11558_/S sky130_fd_sc_hd__buf_4
Xrepeater638 input351/X vssd1 vssd1 vccd1 vccd1 _09185_/C sky130_fd_sc_hd__buf_8
XFILLER_42_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater649 _07986_/A vssd1 vssd1 vccd1 vccd1 _09244_/A sky130_fd_sc_hd__buf_8
XFILLER_38_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06620_ _06620_/A _06620_/B vssd1 vssd1 vccd1 vccd1 _06620_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06551_ _06549_/A _06548_/Y _06549_/Y _06548_/A _06550_/Y vssd1 vssd1 vccd1 vccd1
+ _06552_/B sky130_fd_sc_hd__o221a_1
XFILLER_179_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09270_ _09269_/A _12304_/Q _09268_/B _09269_/X vssd1 vssd1 vccd1 vccd1 _09277_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_61_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06482_ _06522_/A vssd1 vssd1 vccd1 vccd1 _06482_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_61_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08221_ _13082_/Q _08176_/Y _13102_/Q _10460_/A _08220_/X vssd1 vssd1 vccd1 vccd1
+ _08221_/X sky130_fd_sc_hd__o221a_1
XFILLER_53_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08152_ _12831_/Q vssd1 vssd1 vccd1 vccd1 _10477_/A sky130_fd_sc_hd__inv_2
XFILLER_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07103_ _07317_/A _09071_/D _09072_/A _09071_/C vssd1 vssd1 vccd1 vccd1 _09296_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08083_ _08083_/A vssd1 vssd1 vccd1 vccd1 _08083_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07034_ _07046_/A vssd1 vssd1 vccd1 vccd1 _07034_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_173_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13276_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08985_ _09279_/A _09279_/D _09284_/A _08984_/Y vssd1 vssd1 vccd1 vccd1 _08986_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_130_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07936_ _12906_/Q _11495_/X _07946_/S vssd1 vssd1 vccd1 vccd1 _12906_/D sky130_fd_sc_hd__mux2_1
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07867_ _07867_/A _07867_/B _07867_/C _07866_/X vssd1 vssd1 vccd1 vccd1 _07880_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09606_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09611_/A sky130_fd_sc_hd__or2_1
X_06818_ _12019_/X _12018_/X _12019_/X _12018_/X vssd1 vssd1 vccd1 vccd1 _06818_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07798_ _07794_/Y _12923_/Q _07795_/Y _12895_/Q _07797_/X vssd1 vssd1 vccd1 vccd1
+ _07819_/A sky130_fd_sc_hd__a221o_1
XFILLER_83_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09537_ _13176_/Q _13175_/Q _09552_/A _09552_/B vssd1 vssd1 vccd1 vccd1 _09538_/A
+ sky130_fd_sc_hd__o22a_1
X_06749_ _06719_/X _06744_/X _06748_/Y _06480_/X _13203_/Q vssd1 vssd1 vccd1 vccd1
+ _13203_/D sky130_fd_sc_hd__a32o_1
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ _12985_/Q _09436_/X _09008_/B _09451_/X _09467_/X vssd1 vssd1 vccd1 vccd1
+ _09468_/X sky130_fd_sc_hd__a221o_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08419_ _12781_/Q _08417_/X _07997_/X _08418_/X vssd1 vssd1 vccd1 vccd1 _12781_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09399_ _12414_/D vssd1 vssd1 vccd1 vccd1 _09399_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11430_ _12905_/Q _09244_/A _11433_/S vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__mux2_1
XPHY_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11361_ _09327_/A _10533_/Y _12321_/Q vssd1 vssd1 vccd1 vccd1 _11361_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10312_ _10312_/A _11926_/X vssd1 vssd1 vccd1 vccd1 _10312_/Y sky130_fd_sc_hd__nor2b_4
X_13100_ _12167_/X _13100_/D _07236_/X vssd1 vssd1 vccd1 vccd1 _13100_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11292_ vssd1 vssd1 vccd1 vccd1 _11292_/HI _11292_/LO sky130_fd_sc_hd__conb_1
XFILLER_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13031_ _12164_/X _13031_/D _07437_/X vssd1 vssd1 vccd1 vccd1 _13031_/Q sky130_fd_sc_hd__dfrtp_4
X_10243_ _09921_/Y _10134_/X _10234_/X _10242_/X vssd1 vssd1 vccd1 vccd1 _10243_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_65_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10174_ _10045_/A _13146_/Q vssd1 vssd1 vccd1 vccd1 _10174_/X sky130_fd_sc_hd__and2b_1
XFILLER_191_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12815_ _12169_/X _12815_/D _08328_/X vssd1 vssd1 vccd1 vccd1 _12815_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_16_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12746_ _12749_/CLK _12746_/D _08585_/X vssd1 vssd1 vccd1 vccd1 _12746_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _12679_/CLK _12677_/D _08769_/X vssd1 vssd1 vccd1 vccd1 _12677_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11628_ _10498_/X _12927_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11628_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11559_ _12816_/Q _09244_/A _11569_/S vssd1 vssd1 vccd1 vccd1 _11559_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13229_ _13236_/CLK _13229_/D _06487_/X vssd1 vssd1 vccd1 vccd1 _13229_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08770_ _12677_/Q vssd1 vssd1 vccd1 vccd1 _08770_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07721_ _12950_/Q _07717_/X _12949_/Q _07693_/X _07714_/X vssd1 vssd1 vccd1 vccd1
+ _12950_/D sky130_fd_sc_hd__o221a_1
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07652_ _07652_/A _12958_/Q _12959_/Q vssd1 vssd1 vccd1 vccd1 _07652_/X sky130_fd_sc_hd__or3b_1
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06603_ _13219_/Q vssd1 vssd1 vccd1 vccd1 _06603_/Y sky130_fd_sc_hd__inv_2
X_07583_ _08978_/A vssd1 vssd1 vccd1 vccd1 _07583_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09322_ _12367_/Q vssd1 vssd1 vccd1 vccd1 _09330_/A sky130_fd_sc_hd__inv_2
X_06534_ _12761_/Q _12760_/Q vssd1 vssd1 vccd1 vccd1 _06535_/A sky130_fd_sc_hd__and2_1
XFILLER_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09253_ _12456_/Q _09250_/X _10528_/C _09251_/X vssd1 vssd1 vccd1 vccd1 _12456_/D
+ sky130_fd_sc_hd__a22o_1
X_06465_ _06465_/A vssd1 vssd1 vccd1 vccd1 _06465_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08204_ _13088_/Q _10420_/A _08202_/Y _12814_/Q _08203_/X vssd1 vssd1 vccd1 vccd1
+ _08209_/C sky130_fd_sc_hd__a221o_1
X_09184_ _09184_/A _09184_/B vssd1 vssd1 vccd1 vccd1 _09186_/C sky130_fd_sc_hd__or2_1
XFILLER_166_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06396_ _06396_/A vssd1 vssd1 vccd1 vccd1 _06396_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08135_ _12814_/Q vssd1 vssd1 vccd1 vccd1 _10433_/B sky130_fd_sc_hd__inv_2
XFILLER_162_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08066_ _08082_/A vssd1 vssd1 vccd1 vccd1 _08066_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07017_ _06886_/X _12185_/X _06887_/X _13169_/Q vssd1 vssd1 vccd1 vccd1 _13169_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput205 la_oenb[19] vssd1 vssd1 vccd1 vccd1 input205/X sky130_fd_sc_hd__buf_1
Xinput216 la_oenb[29] vssd1 vssd1 vccd1 vccd1 input216/X sky130_fd_sc_hd__buf_1
Xinput227 la_oenb[39] vssd1 vssd1 vccd1 vccd1 input227/X sky130_fd_sc_hd__buf_1
Xinput238 la_oenb[49] vssd1 vssd1 vccd1 vccd1 input238/X sky130_fd_sc_hd__buf_1
X_08968_ _08969_/A vssd1 vssd1 vccd1 vccd1 _08968_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput249 la_oenb[59] vssd1 vssd1 vccd1 vccd1 input249/X sky130_fd_sc_hd__buf_1
XFILLER_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07919_ _07933_/A vssd1 vssd1 vccd1 vccd1 _07931_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08899_ _08898_/X _06316_/A _08893_/X _12629_/Q vssd1 vssd1 vccd1 vccd1 _12629_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_112_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10930_ _10930_/A _10930_/B vssd1 vssd1 vccd1 vccd1 _10930_/Y sky130_fd_sc_hd__nor2_4
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_92_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _13156_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_21_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12619_/CLK sky130_fd_sc_hd__clkbuf_16
X_10861_ _12522_/Q vssd1 vssd1 vccd1 vccd1 _10861_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12600_ _12975_/CLK _12600_/D vssd1 vssd1 vccd1 vccd1 _12600_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ _10792_/A _10792_/B _10792_/C _10792_/D vssd1 vssd1 vccd1 vccd1 _10796_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_52_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12537_/CLK _12531_/D vssd1 vssd1 vccd1 vccd1 _12531_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12462_ _12985_/CLK _12462_/D vssd1 vssd1 vccd1 vccd1 _12462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11413_ _11412_/X _12443_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11413_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12393_ _12413_/CLK _12393_/D vssd1 vssd1 vccd1 vccd1 _12415_/D sky130_fd_sc_hd__dfxtp_2
X_11344_ _11344_/A vssd1 vssd1 vccd1 vccd1 _11344_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ vssd1 vssd1 vccd1 vccd1 _11275_/HI _11275_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13014_ _12164_/X _13014_/D _07481_/X vssd1 vssd1 vccd1 vccd1 _13014_/Q sky130_fd_sc_hd__dfrtp_4
X_10226_ _10214_/Y _10134_/X _10217_/X _10225_/X vssd1 vssd1 vccd1 vccd1 _10226_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10157_ _13261_/Q vssd1 vssd1 vccd1 vccd1 _10157_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10088_ _10088_/A _10088_/B _10088_/C _10088_/D vssd1 vssd1 vccd1 vccd1 _10088_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12729_ _12735_/CLK _12729_/D _08630_/X vssd1 vssd1 vccd1 vccd1 _12729_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06250_ _08996_/D vssd1 vssd1 vccd1 vccd1 _06280_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06181_ _06092_/A _06132_/B _06179_/Y _06077_/Y _06180_/X vssd1 vssd1 vccd1 vccd1
+ _06181_/X sky130_fd_sc_hd__o311a_2
XFILLER_144_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09940_ _09950_/A vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__clkbuf_2
X_09871_ _09879_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _09877_/A sky130_fd_sc_hd__or2_1
XFILLER_48_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08822_ _08814_/X _08817_/X _06323_/Y _12660_/Q _08811_/X vssd1 vssd1 vccd1 vccd1
+ _12660_/D sky130_fd_sc_hd__a32o_1
XFILLER_86_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08753_ _12682_/Q vssd1 vssd1 vccd1 vccd1 _08753_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07704_ _12959_/Q _07694_/X _07698_/X _07702_/Y _07703_/X vssd1 vssd1 vccd1 vccd1
+ _12959_/D sky130_fd_sc_hd__o221a_1
XPHY_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08684_/X sky130_fd_sc_hd__buf_1
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07635_ _12954_/Q vssd1 vssd1 vccd1 vccd1 _07665_/B sky130_fd_sc_hd__inv_2
XPHY_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07566_ _09226_/B vssd1 vssd1 vccd1 vccd1 _07566_/X sky130_fd_sc_hd__buf_4
XFILLER_22_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09305_ _08877_/X _07737_/X _07732_/X _12618_/Q _07037_/X vssd1 vssd1 vccd1 vccd1
+ _12618_/D sky130_fd_sc_hd__a41o_1
X_06517_ _06517_/A vssd1 vssd1 vccd1 vccd1 _06527_/A sky130_fd_sc_hd__inv_2
XFILLER_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07497_ _11982_/X vssd1 vssd1 vccd1 vccd1 _07497_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09236_ _12464_/Q _09233_/A _07558_/X _09083_/X vssd1 vssd1 vccd1 vccd1 _12464_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06448_ _12116_/X vssd1 vssd1 vccd1 vccd1 _06448_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09167_ _11626_/X _09163_/X _12501_/Q _09164_/X vssd1 vssd1 vccd1 vccd1 _12501_/D
+ sky130_fd_sc_hd__a22o_1
X_06379_ _13248_/Q vssd1 vssd1 vccd1 vccd1 _06379_/X sky130_fd_sc_hd__buf_2
XFILLER_5_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08118_ _08114_/Y _10475_/A _08116_/Y _08117_/X vssd1 vssd1 vccd1 vccd1 _08118_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09098_ _12536_/Q _09089_/X _10794_/D _09092_/X vssd1 vssd1 vccd1 vccd1 _12536_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08049_ _08051_/A vssd1 vssd1 vccd1 vccd1 _08049_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_150_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11060_ _11899_/X vssd1 vssd1 vccd1 vccd1 _11060_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10011_ _08748_/Y _10134_/A _06191_/Y _09972_/A _09991_/A vssd1 vssd1 vccd1 vccd1
+ _10011_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_103_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11962_ _07746_/X _09259_/Y _12607_/Q vssd1 vssd1 vccd1 vccd1 _11962_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10913_ _12529_/Q _12341_/Q _10911_/Y _10912_/Y vssd1 vssd1 vccd1 vccd1 _10915_/A
+ sky130_fd_sc_hd__o22a_2
X_11893_ _10775_/X _10753_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _11893_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ _10843_/A _10843_/B _10843_/Y vssd1 vssd1 vccd1 vccd1 _10847_/A sky130_fd_sc_hd__a21oi_2
XFILLER_13_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10775_ _10736_/X _10750_/X _06365_/X _10751_/X _10752_/X vssd1 vssd1 vccd1 vccd1
+ _10775_/X sky130_fd_sc_hd__a221o_1
XFILLER_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12514_ _12849_/CLK _12514_/D vssd1 vssd1 vccd1 vccd1 _12514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12445_ _12489_/CLK _12445_/D vssd1 vssd1 vccd1 vccd1 _12445_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12376_ _12376_/CLK _12376_/D vssd1 vssd1 vccd1 vccd1 _12398_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_158_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput509 _11257_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11327_ vssd1 vssd1 vccd1 vccd1 _11327_/HI _11327_/LO sky130_fd_sc_hd__conb_1
XFILLER_114_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11258_ vssd1 vssd1 vccd1 vccd1 _11258_/HI _11258_/LO sky130_fd_sc_hd__conb_1
XFILLER_140_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10209_ _10208_/Y _10045_/A _08159_/Y _10113_/X vssd1 vssd1 vccd1 vccd1 _10209_/X
+ sky130_fd_sc_hd__o22a_1
X_11189_ vssd1 vssd1 vccd1 vccd1 _11189_/HI _11189_/LO sky130_fd_sc_hd__conb_1
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07420_ _07428_/A vssd1 vssd1 vccd1 vccd1 _07420_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07351_ _11438_/X _07338_/X _13062_/Q _07339_/X vssd1 vssd1 vccd1 vccd1 _13062_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06302_ _06313_/A vssd1 vssd1 vccd1 vccd1 _06302_/X sky130_fd_sc_hd__clkbuf_1
X_07282_ _07362_/A vssd1 vssd1 vccd1 vccd1 _07302_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_176_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09021_ _09023_/A input38/X vssd1 vssd1 vccd1 vccd1 _12577_/D sky130_fd_sc_hd__and2_1
X_06233_ _06050_/X _06232_/Y _06050_/X _06232_/Y vssd1 vssd1 vccd1 vccd1 _06233_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_191_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06164_ _06005_/Y _06022_/X _11963_/S _06163_/X vssd1 vssd1 vccd1 vccd1 _13286_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_172_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06095_ _12728_/Q _12696_/Q _12727_/Q _12695_/Q vssd1 vssd1 vccd1 vccd1 _06095_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09923_ _12887_/Q _09935_/B vssd1 vssd1 vccd1 vccd1 _09923_/X sky130_fd_sc_hd__or2_1
XFILLER_160_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09854_ _09866_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09860_/A sky130_fd_sc_hd__or2_1
XFILLER_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08805_ _08807_/A vssd1 vssd1 vccd1 vccd1 _08805_/X sky130_fd_sc_hd__clkbuf_1
X_09785_ _09785_/A _09802_/A vssd1 vssd1 vccd1 vccd1 _09785_/X sky130_fd_sc_hd__or2_1
XFILLER_74_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06997_ _07006_/A vssd1 vssd1 vccd1 vccd1 _06997_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08736_ _08747_/A vssd1 vssd1 vccd1 vccd1 _08736_/X sky130_fd_sc_hd__clkbuf_1
XPHY_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _08669_/A vssd1 vssd1 vccd1 vccd1 _08667_/X sky130_fd_sc_hd__clkbuf_1
XPHY_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07618_ _11613_/X _07610_/X _12968_/Q _07611_/X _07616_/X vssd1 vssd1 vccd1 vccd1
+ _12968_/D sky130_fd_sc_hd__o221a_1
XPHY_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _08606_/A vssd1 vssd1 vccd1 vccd1 _08598_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ _07549_/A vssd1 vssd1 vccd1 vccd1 _11356_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_139_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10560_ _10608_/A _10608_/B vssd1 vssd1 vccd1 vccd1 _11392_/S sky130_fd_sc_hd__or2_4
XFILLER_128_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ _12472_/Q _09215_/X _07562_/X _09216_/X vssd1 vssd1 vccd1 vccd1 _12472_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10491_ _12496_/Q _09135_/B _09136_/B vssd1 vssd1 vccd1 vccd1 _10491_/X sky130_fd_sc_hd__a21bo_1
XFILLER_5_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12230_ _12229_/X _12635_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12230_/X sky130_fd_sc_hd__mux2_2
XFILLER_108_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12161_ _10786_/X _11143_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _12161_/X sky130_fd_sc_hd__mux2_2
XFILLER_150_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11112_ _12116_/X vssd1 vssd1 vccd1 vccd1 _11112_/X sky130_fd_sc_hd__clkbuf_2
X_12092_ _12448_/Q _12091_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _12092_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11043_ _10699_/X _11037_/X _06400_/X _07020_/X _11038_/X vssd1 vssd1 vccd1 vccd1
+ _11043_/X sky130_fd_sc_hd__a221o_1
XFILLER_89_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12994_ _12999_/CLK _12994_/D vssd1 vssd1 vccd1 vccd1 _12994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11945_ _09735_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11945_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11876_ _10293_/X _12817_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11876_/X sky130_fd_sc_hd__mux2_2
XFILLER_44_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10827_ _10827_/A vssd1 vssd1 vccd1 vccd1 _10827_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10758_ _10758_/A vssd1 vssd1 vccd1 vccd1 _10758_/X sky130_fd_sc_hd__buf_2
XFILLER_185_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10689_ _10701_/A _10691_/B _10688_/X vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__o21a_1
XFILLER_195_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12428_ _12471_/CLK _12428_/D vssd1 vssd1 vccd1 vccd1 _12428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12359_ _13257_/CLK _12359_/D vssd1 vssd1 vccd1 vccd1 _12359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06920_ _07026_/A vssd1 vssd1 vccd1 vccd1 _06973_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06851_ _06848_/X _06849_/X _12030_/X _06850_/X vssd1 vssd1 vccd1 vccd1 _06851_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09570_ _09569_/Y _07735_/A _12869_/Q _07729_/X vssd1 vssd1 vccd1 vccd1 _09570_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06782_ _12008_/X _06751_/X _12008_/X _06751_/X vssd1 vssd1 vccd1 vccd1 _06783_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_08521_ _08521_/A vssd1 vssd1 vccd1 vccd1 _08533_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_149_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12802_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08452_ _13048_/Q _10333_/A _08450_/Y _12903_/Q _08451_/X vssd1 vssd1 vccd1 vccd1
+ _08457_/C sky130_fd_sc_hd__a221o_1
XFILLER_1_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07403_ _12841_/Q vssd1 vssd1 vccd1 vccd1 _07403_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08383_ _08385_/A vssd1 vssd1 vccd1 vccd1 _08383_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_189_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07334_ _11445_/X _07321_/X _13069_/Q _07324_/X vssd1 vssd1 vccd1 vccd1 _13069_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07265_ _11554_/X _07263_/X _13089_/Q _07264_/X vssd1 vssd1 vccd1 vccd1 _13089_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09004_ _09008_/A _09008_/B _11648_/X vssd1 vssd1 vccd1 vccd1 _12592_/D sky130_fd_sc_hd__and3_1
XFILLER_136_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06216_ _06281_/A vssd1 vssd1 vccd1 vccd1 _06216_/X sky130_fd_sc_hd__clkbuf_2
X_07196_ _09984_/A _09982_/B _09302_/A vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__or3_4
XFILLER_117_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06147_ _12742_/Q _12710_/Q _06146_/X vssd1 vssd1 vccd1 vccd1 _06147_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_118_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06078_ _12732_/Q _12700_/Q _12731_/Q _12699_/Q vssd1 vssd1 vccd1 vccd1 _06078_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09906_ _12659_/Q vssd1 vssd1 vccd1 vccd1 _09906_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09837_ _09837_/A vssd1 vssd1 vccd1 vccd1 _09837_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09768_ _09886_/A _09768_/B vssd1 vssd1 vccd1 vccd1 _09768_/X sky130_fd_sc_hd__or2_1
XFILLER_74_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _08729_/A vssd1 vssd1 vccd1 vccd1 _08719_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_199_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09699_ _09713_/B _09698_/Y _09696_/A _09698_/A _09701_/A vssd1 vssd1 vccd1 vccd1
+ _09700_/B sky130_fd_sc_hd__o221a_1
XFILLER_199_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11729_/X _11922_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12442_/D sky130_fd_sc_hd__mux2_1
XPHY_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11384_/X _09184_/A _11675_/S vssd1 vssd1 vccd1 vccd1 _11661_/X sky130_fd_sc_hd__mux2_1
XPHY_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10612_ _10612_/A vssd1 vssd1 vccd1 vccd1 _10619_/B sky130_fd_sc_hd__buf_1
XFILLER_70_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ _10442_/Y _10528_/C _11592_/S vssd1 vssd1 vccd1 vccd1 _11592_/X sky130_fd_sc_hd__mux2_1
XPHY_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10543_ _11359_/X vssd1 vssd1 vccd1 vccd1 _10543_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13262_ _13264_/CLK _13262_/D _06313_/X vssd1 vssd1 vccd1 vccd1 _13262_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10474_ _10474_/A _10475_/B _10474_/C vssd1 vssd1 vccd1 vccd1 _10474_/Y sky130_fd_sc_hd__nor3_1
XFILLER_182_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12213_ _06327_/Y _13152_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12213_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13193_ _13193_/CLK _13193_/D _06839_/X vssd1 vssd1 vccd1 vccd1 _13193_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ _09992_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _12144_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12075_ _12446_/Q _12074_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _12075_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11026_ _07888_/Y _08494_/X _12841_/Q vssd1 vssd1 vccd1 vccd1 _12551_/D sky130_fd_sc_hd__o21a_1
XFILLER_92_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12977_ _12977_/CLK _12977_/D vssd1 vssd1 vccd1 vccd1 _12977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11928_ _09486_/X _12789_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11928_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11859_ _10092_/Y _12806_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11859_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07050_ _07063_/A vssd1 vssd1 vccd1 vccd1 _07050_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07952_ _07804_/X _11489_/X _07962_/S vssd1 vssd1 vccd1 vccd1 _12900_/D sky130_fd_sc_hd__mux2_1
XFILLER_87_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06903_ _06900_/X _06901_/X _12028_/X _06902_/X vssd1 vssd1 vccd1 vccd1 _06903_/X
+ sky130_fd_sc_hd__o22a_1
X_07883_ _09302_/A _09981_/C vssd1 vssd1 vccd1 vccd1 _09969_/B sky130_fd_sc_hd__or2_4
XFILLER_56_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09622_ _09614_/Y _09621_/Y _09614_/Y _09621_/Y vssd1 vssd1 vccd1 vccd1 _09625_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_06834_ _12031_/X _06840_/B vssd1 vssd1 vccd1 vccd1 _06834_/X sky130_fd_sc_hd__or2_2
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09553_ _09552_/A _09552_/B _09552_/C vssd1 vssd1 vccd1 vccd1 _09554_/B sky130_fd_sc_hd__o21a_1
XFILLER_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06765_ _06765_/A vssd1 vssd1 vccd1 vccd1 _13202_/D sky130_fd_sc_hd__inv_2
XFILLER_71_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08504_ _08504_/A vssd1 vssd1 vccd1 vccd1 _08504_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09484_ _13148_/Q vssd1 vssd1 vccd1 vccd1 _09484_/Y sky130_fd_sc_hd__inv_2
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06696_ _11034_/A vssd1 vssd1 vccd1 vccd1 _10687_/A sky130_fd_sc_hd__inv_2
XFILLER_52_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08435_ _08521_/A vssd1 vssd1 vccd1 vccd1 _08503_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ _08370_/A vssd1 vssd1 vccd1 vccd1 _08366_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_149_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07317_ _07317_/A _09042_/B vssd1 vssd1 vccd1 vccd1 _09295_/A sky130_fd_sc_hd__or2_4
XFILLER_176_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08297_ _12828_/Q _11603_/X _08307_/S vssd1 vssd1 vccd1 vccd1 _12828_/D sky130_fd_sc_hd__mux2_1
XFILLER_164_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07248_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07248_/X sky130_fd_sc_hd__buf_2
XFILLER_125_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12464_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07179_ _07183_/A vssd1 vssd1 vccd1 vccd1 _07179_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_127_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10190_ _10190_/A _11979_/X vssd1 vssd1 vccd1 vccd1 _10190_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_133_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12900_ _12166_/X _12900_/D _07950_/X vssd1 vssd1 vccd1 vccd1 _12900_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12831_ _12169_/X _12831_/D _08289_/X vssd1 vssd1 vccd1 vccd1 _12831_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12762_ _12779_/CLK _12762_/D _08516_/X vssd1 vssd1 vccd1 vccd1 _12762_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_199_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11713_ _10641_/Y _10642_/Y _11818_/S vssd1 vssd1 vccd1 vccd1 _11713_/X sky130_fd_sc_hd__mux2_1
XPHY_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12693_ _12725_/CLK _12693_/D _08721_/X vssd1 vssd1 vccd1 vccd1 _12693_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_187_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _10514_/X _12929_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11644_/X sky130_fd_sc_hd__mux2_1
XPHY_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 io_in[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_1
XFILLER_7_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11575_ _12832_/Q _10794_/B _11578_/S vssd1 vssd1 vccd1 vccd1 _11575_/X sky130_fd_sc_hd__mux2_1
Xinput27 io_in[33] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_1
XFILLER_11_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput38 io_in[9] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_1
XFILLER_196_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10526_ _10526_/A _10526_/B vssd1 vssd1 vccd1 vccd1 _10526_/Y sky130_fd_sc_hd__nor2_1
Xinput49 la_data_in[109] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_1
XFILLER_109_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13245_ _13249_/CLK _13245_/D _06388_/X vssd1 vssd1 vccd1 vccd1 _13245_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_7_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10457_ _10454_/B _10450_/A _10454_/A vssd1 vssd1 vccd1 vccd1 _10458_/C sky130_fd_sc_hd__o21a_1
XFILLER_108_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13176_ _13177_/CLK _13176_/D _06981_/X vssd1 vssd1 vccd1 vccd1 _13176_/Q sky130_fd_sc_hd__dfrtp_4
X_10388_ _10388_/A _10388_/B vssd1 vssd1 vccd1 vccd1 _10390_/B sky130_fd_sc_hd__nand2_2
XFILLER_123_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12127_ _12126_/X _12437_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12127_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12058_ _12439_/Q _12057_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12058_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater617 _11492_/S vssd1 vssd1 vccd1 vccd1 _11501_/S sky130_fd_sc_hd__buf_4
XFILLER_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater628 _11543_/S vssd1 vssd1 vccd1 vccd1 _11533_/S sky130_fd_sc_hd__buf_6
Xrepeater639 input342/X vssd1 vssd1 vccd1 vccd1 _09180_/A sky130_fd_sc_hd__buf_8
X_11009_ _12356_/Q vssd1 vssd1 vccd1 vccd1 _11013_/A sky130_fd_sc_hd__inv_2
XFILLER_133_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06550_ _06540_/X _06544_/X _06552_/A vssd1 vssd1 vccd1 vccd1 _06550_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_179_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06481_ _06457_/X _06473_/X _06479_/Y _06480_/X _13231_/Q vssd1 vssd1 vccd1 vccd1
+ _13231_/D sky130_fd_sc_hd__a32o_1
XFILLER_61_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08220_ _13094_/Q _08187_/X _13094_/Q _08187_/X vssd1 vssd1 vccd1 vccd1 _08220_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_178_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08151_ _08151_/A _08151_/B _08151_/C _08150_/X vssd1 vssd1 vccd1 vccd1 _08163_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_119_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07102_ _07102_/A _07102_/B _07102_/C _07102_/D vssd1 vssd1 vccd1 vccd1 _09072_/A
+ sky130_fd_sc_hd__or4_4
X_08082_ _08082_/A vssd1 vssd1 vccd1 vccd1 _08082_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07033_ _06663_/X _12182_/X _06415_/B _13163_/Q vssd1 vssd1 vccd1 vccd1 _13163_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_146_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08984_ _12304_/Q vssd1 vssd1 vccd1 vccd1 _08984_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07935_ _07967_/S vssd1 vssd1 vccd1 vccd1 _07946_/S sky130_fd_sc_hd__buf_2
XFILLER_60_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_164_wb_clk_i clkbuf_opt_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _12558_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07866_ _07859_/X _07866_/B _07866_/C _07866_/D vssd1 vssd1 vccd1 vccd1 _07866_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_113_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09605_ _09604_/A _09604_/B _09604_/C vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__o21a_1
X_06817_ _12010_/X _06815_/B _06815_/X vssd1 vssd1 vccd1 vccd1 _06817_/X sky130_fd_sc_hd__a21bo_1
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07797_ _13013_/Q _10328_/A _13013_/Q _10328_/A vssd1 vssd1 vccd1 vccd1 _07797_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09536_ _13176_/Q vssd1 vssd1 vccd1 vccd1 _09552_/A sky130_fd_sc_hd__inv_2
X_06748_ _06748_/A _06748_/B vssd1 vssd1 vccd1 vccd1 _06748_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ _12973_/Q _09440_/X _12933_/Q _09438_/A _09466_/X vssd1 vssd1 vccd1 vccd1
+ _09467_/X sky130_fd_sc_hd__a221o_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06679_ _06672_/Y _12051_/X _06673_/X _06680_/A vssd1 vssd1 vccd1 vccd1 _06679_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08418_ _08418_/A vssd1 vssd1 vccd1 vccd1 _08418_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_197_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09398_ _12398_/D vssd1 vssd1 vccd1 vccd1 _10562_/A sky130_fd_sc_hd__inv_2
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08349_ _12806_/Q _11581_/X _08349_/S vssd1 vssd1 vccd1 vccd1 _12806_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11360_ _09328_/A _10538_/X _12321_/Q vssd1 vssd1 vccd1 vccd1 _11360_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10311_ _10310_/Y _09972_/A _09937_/Y _09968_/X _09991_/A vssd1 vssd1 vccd1 vccd1
+ _10311_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_152_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11291_ vssd1 vssd1 vccd1 vccd1 _11291_/HI _11291_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13030_ _12164_/X _13030_/D _07439_/X vssd1 vssd1 vccd1 vccd1 _13030_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10242_ _10235_/Y _10140_/X _10236_/Y _10141_/X _10241_/X vssd1 vssd1 vccd1 vccd1
+ _10242_/X sky130_fd_sc_hd__o221a_1
XFILLER_152_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10173_ _10190_/A _11978_/X vssd1 vssd1 vccd1 vccd1 _10173_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_154_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12814_ _12169_/X _12814_/D _08330_/X vssd1 vssd1 vccd1 vccd1 _12814_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_43_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12745_ _12747_/CLK _12745_/D _08587_/X vssd1 vssd1 vccd1 vccd1 _12745_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_43_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12679_/CLK _12676_/D _08773_/X vssd1 vssd1 vccd1 vccd1 _12676_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_169_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _10497_/X _12926_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11627_/X sky130_fd_sc_hd__mux2_1
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ _12815_/Q _09244_/B _11558_/S vssd1 vssd1 vccd1 vccd1 _11558_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10509_ _12583_/Q _07757_/B _07758_/B vssd1 vssd1 vccd1 vccd1 _10509_/X sky130_fd_sc_hd__a21bo_1
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11489_ _10336_/X input358/X _11492_/S vssd1 vssd1 vccd1 vccd1 _11489_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13228_ _13237_/CLK _13228_/D _06502_/X vssd1 vssd1 vccd1 vccd1 _13228_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13159_ _13159_/CLK _13159_/D _07050_/X vssd1 vssd1 vccd1 vccd1 _13159_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07720_ _12951_/Q _07717_/X _07698_/X _07719_/Y _07714_/X vssd1 vssd1 vccd1 vccd1
+ _12951_/D sky130_fd_sc_hd__o221a_1
XFILLER_84_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07651_ _12951_/Q _07651_/B _12950_/Q vssd1 vssd1 vccd1 vccd1 _08980_/A sky130_fd_sc_hd__or3b_4
XFILLER_93_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_168_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06602_ _06602_/A _06602_/B vssd1 vssd1 vccd1 vccd1 _06602_/Y sky130_fd_sc_hd__nor2_1
X_07582_ _12980_/Q _07574_/X _09226_/A _07575_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _12980_/D sky130_fd_sc_hd__o221a_1
X_09321_ _12368_/Q vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__inv_2
X_06533_ _13224_/Q vssd1 vssd1 vccd1 vccd1 _06533_/Y sky130_fd_sc_hd__inv_2
X_09252_ _12457_/Q _09250_/X _09243_/A _09251_/X vssd1 vssd1 vccd1 vccd1 _12457_/D
+ sky130_fd_sc_hd__a22o_1
X_06464_ _06440_/X _06462_/Y _06420_/X _06463_/Y vssd1 vssd1 vccd1 vccd1 _13233_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_194_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08203_ _13113_/Q _08122_/Y _13095_/Q _10439_/A vssd1 vssd1 vccd1 vccd1 _08203_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09183_ _09183_/A _10528_/B _10529_/A _09183_/D vssd1 vssd1 vccd1 vccd1 _09187_/C
+ sky130_fd_sc_hd__or4_4
X_06395_ _06412_/A vssd1 vssd1 vccd1 vccd1 _06395_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_159_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08134_ _13136_/Q _10467_/B _13074_/Q vssd1 vssd1 vccd1 vccd1 _08163_/A sky130_fd_sc_hd__o21ai_1
XFILLER_119_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08065_ _08067_/A vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__buf_2
XFILLER_174_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07016_ _07024_/A vssd1 vssd1 vccd1 vccd1 _07016_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_89_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput206 la_oenb[1] vssd1 vssd1 vccd1 vccd1 _11345_/A sky130_fd_sc_hd__buf_4
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput217 la_oenb[2] vssd1 vssd1 vccd1 vccd1 input217/X sky130_fd_sc_hd__buf_1
XFILLER_103_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput228 la_oenb[3] vssd1 vssd1 vccd1 vccd1 input228/X sky130_fd_sc_hd__buf_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08967_ _08969_/A vssd1 vssd1 vccd1 vccd1 _08967_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput239 la_oenb[4] vssd1 vssd1 vccd1 vccd1 input239/X sky130_fd_sc_hd__buf_1
X_07918_ _12913_/Q _11502_/X _07918_/S vssd1 vssd1 vccd1 vccd1 _12913_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08898_ _08898_/A vssd1 vssd1 vccd1 vccd1 _08898_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07849_ _13019_/Q _10346_/B _13014_/Q _10331_/A _07848_/X vssd1 vssd1 vccd1 vccd1
+ _07867_/B sky130_fd_sc_hd__a221o_1
XFILLER_56_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10860_ _10858_/A _10859_/A _10864_/C _10859_/Y vssd1 vssd1 vccd1 vccd1 _12333_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_83_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09519_ _09510_/Y _07069_/A _12865_/Q _07729_/X _09518_/X vssd1 vssd1 vccd1 vccd1
+ _09519_/X sky130_fd_sc_hd__a221o_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _10755_/X _10737_/X _06371_/X _10738_/X _10739_/X vssd1 vssd1 vccd1 vccd1
+ _10791_/X sky130_fd_sc_hd__a221o_1
XFILLER_140_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12537_/CLK _12530_/D vssd1 vssd1 vccd1 vccd1 _12530_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_wb_clk_i _12960_/CLK vssd1 vssd1 vccd1 vccd1 _13243_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _12464_/CLK _12461_/D vssd1 vssd1 vccd1 vccd1 _12461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11412_ _12443_/Q _11411_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _11412_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12392_ _12995_/CLK _12392_/D vssd1 vssd1 vccd1 vccd1 _12414_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11343_ vssd1 vssd1 vccd1 vccd1 _11343_/HI _11343_/LO sky130_fd_sc_hd__conb_1
XFILLER_67_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11274_ vssd1 vssd1 vccd1 vccd1 _11274_/HI _11274_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13013_ _12164_/X _13013_/D _07483_/X vssd1 vssd1 vccd1 vccd1 _13013_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10225_ _10218_/Y _10140_/X _09584_/Y _10141_/X _10224_/X vssd1 vssd1 vccd1 vccd1
+ _10225_/X sky130_fd_sc_hd__o221a_1
XFILLER_152_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10156_ _10015_/B _08984_/Y _09279_/B _09279_/X vssd1 vssd1 vccd1 vccd1 _12304_/D
+ sky130_fd_sc_hd__o31ai_1
XFILLER_43_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10087_ _10083_/Y _09999_/A _09494_/Y _10141_/A _10086_/X vssd1 vssd1 vccd1 vccd1
+ _10088_/D sky130_fd_sc_hd__o221a_1
XFILLER_75_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10989_ _12538_/Q _12350_/Q _12539_/Q _12351_/Q vssd1 vssd1 vccd1 vccd1 _10989_/X
+ sky130_fd_sc_hd__a22o_1
X_12728_ _12735_/CLK _12728_/D _08632_/X vssd1 vssd1 vccd1 vccd1 _12728_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12659_ _12664_/CLK _12659_/D _08823_/X vssd1 vssd1 vccd1 vccd1 _12659_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06180_ _06180_/A _06180_/B _06096_/X vssd1 vssd1 vccd1 vccd1 _06180_/X sky130_fd_sc_hd__or3b_2
XFILLER_117_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09870_ _09879_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _09870_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08821_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08821_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08752_ _08769_/A vssd1 vssd1 vccd1 vccd1 _08752_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07703_ _09268_/B vssd1 vssd1 vccd1 vccd1 _07703_/X sky130_fd_sc_hd__buf_2
X_08683_ _11842_/X _08670_/X _12708_/Q _08671_/X vssd1 vssd1 vccd1 vccd1 _12708_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07634_ _12962_/Q _07660_/D vssd1 vssd1 vccd1 vccd1 _07646_/D sky130_fd_sc_hd__or2_2
XFILLER_93_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07565_ _07564_/X _07552_/X _12988_/Q _07553_/X _07556_/X vssd1 vssd1 vccd1 vccd1
+ _12988_/D sky130_fd_sc_hd__a221o_1
XFILLER_59_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09304_ _09304_/A _09304_/B vssd1 vssd1 vccd1 vccd1 _11803_/S sky130_fd_sc_hd__nor2_2
XFILLER_0_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06516_ _12162_/X _12161_/X _12160_/X _11959_/X _06520_/A vssd1 vssd1 vccd1 vccd1
+ _06517_/A sky130_fd_sc_hd__a41o_1
XFILLER_22_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07496_ _09185_/A vssd1 vssd1 vccd1 vccd1 _09228_/A sky130_fd_sc_hd__inv_2
XFILLER_55_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09235_ _12465_/Q _09231_/X _07536_/X _09233_/X vssd1 vssd1 vccd1 vccd1 _12465_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06447_ _10711_/A vssd1 vssd1 vccd1 vccd1 _06860_/A sky130_fd_sc_hd__inv_2
XFILLER_166_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09166_ _11627_/X _09163_/X _12502_/Q _09164_/X vssd1 vssd1 vccd1 vccd1 _12502_/D
+ sky130_fd_sc_hd__a22o_1
X_06378_ _06391_/A vssd1 vssd1 vccd1 vccd1 _06378_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_148_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08117_ _12811_/Q vssd1 vssd1 vccd1 vccd1 _08117_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09097_ _12537_/Q _09089_/X _10794_/C _09092_/X vssd1 vssd1 vccd1 vccd1 _12537_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08048_ _12867_/Q _08040_/X _08005_/X _08041_/X vssd1 vssd1 vccd1 vccd1 _12867_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10010_ _10010_/A vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__buf_2
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09999_ _09999_/A vssd1 vssd1 vccd1 vccd1 _10000_/A sky130_fd_sc_hd__buf_2
XFILLER_130_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11961_ _08740_/A _09259_/Y _12607_/Q vssd1 vssd1 vccd1 vccd1 _11961_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10912_ _12341_/Q vssd1 vssd1 vccd1 vccd1 _10912_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11892_ _10776_/X _10762_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _11892_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10843_ _10843_/A _10843_/B vssd1 vssd1 vccd1 vccd1 _10843_/Y sky130_fd_sc_hd__nor2_2
XFILLER_198_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10774_ _10773_/X _10768_/X _06386_/X _10769_/X _10770_/X vssd1 vssd1 vccd1 vccd1
+ _10774_/X sky130_fd_sc_hd__a221o_1
XFILLER_34_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12513_ _12999_/CLK _12513_/D vssd1 vssd1 vccd1 vccd1 _12513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12444_ _12489_/CLK _12444_/D vssd1 vssd1 vccd1 vccd1 _12444_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12375_ _12415_/CLK _12375_/D vssd1 vssd1 vccd1 vccd1 _12397_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11326_ vssd1 vssd1 vccd1 vccd1 _11326_/HI _11326_/LO sky130_fd_sc_hd__conb_1
XFILLER_5_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11257_ vssd1 vssd1 vccd1 vccd1 _11257_/HI _11257_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10208_ hold1/A vssd1 vssd1 vccd1 vccd1 _10208_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11188_ vssd1 vssd1 vccd1 vccd1 _11188_/HI _11188_/LO sky130_fd_sc_hd__conb_1
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10139_ _12777_/Q vssd1 vssd1 vccd1 vccd1 _10139_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07350_ _07360_/A vssd1 vssd1 vccd1 vccd1 _07350_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06301_ _06269_/X _06281_/X _06300_/Y _13265_/Q _06273_/X vssd1 vssd1 vccd1 vccd1
+ _13265_/D sky130_fd_sc_hd__a32o_1
XFILLER_149_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07281_ _11547_/X _07248_/A _13082_/Q _07249_/A vssd1 vssd1 vccd1 vccd1 _13082_/D
+ sky130_fd_sc_hd__a22o_1
X_09020_ _09023_/A _12577_/Q vssd1 vssd1 vccd1 vccd1 _12578_/D sky130_fd_sc_hd__and2_1
XFILLER_148_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06232_ _06047_/Y _06048_/Y _06051_/A _06184_/X vssd1 vssd1 vccd1 vccd1 _06232_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_191_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06163_ _06217_/A vssd1 vssd1 vccd1 vccd1 _06163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06094_ _12726_/Q _12694_/Q _06093_/X vssd1 vssd1 vccd1 vccd1 _06094_/X sky130_fd_sc_hd__o21a_1
XFILLER_172_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09922_ _09952_/A vssd1 vssd1 vccd1 vccd1 _09922_/X sky130_fd_sc_hd__clkbuf_2
X_09853_ _09866_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09853_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08804_ _08798_/X _08801_/X _06283_/Y _12667_/Q _08567_/X vssd1 vssd1 vccd1 vccd1
+ _12667_/D sky130_fd_sc_hd__a32o_1
XFILLER_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09784_ _09785_/A _09802_/A vssd1 vssd1 vccd1 vccd1 _09784_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06996_ _06528_/X _06991_/Y _06995_/X _06841_/X _13174_/Q vssd1 vssd1 vccd1 vccd1
+ _13174_/D sky130_fd_sc_hd__a32o_1
XFILLER_105_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08735_ _11821_/X _08592_/A _12687_/Q _08593_/A vssd1 vssd1 vccd1 vccd1 _12687_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _11849_/X _08654_/X _12715_/Q _08655_/X vssd1 vssd1 vccd1 vccd1 _12715_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07617_ _11614_/X _07610_/X _12969_/Q _07611_/X _07616_/X vssd1 vssd1 vccd1 vccd1
+ _12969_/D sky130_fd_sc_hd__o221a_1
XPHY_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08597_ _11951_/X _08592_/X _12742_/Q _08593_/X vssd1 vssd1 vccd1 vccd1 _12742_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07548_ _09441_/A _09435_/B _09986_/B vssd1 vssd1 vccd1 vccd1 _07549_/A sky130_fd_sc_hd__and3_1
XPHY_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07479_ _07489_/A vssd1 vssd1 vccd1 vccd1 _07479_/X sky130_fd_sc_hd__clkbuf_1
X_09218_ _12473_/Q _09215_/X _07560_/X _09216_/X vssd1 vssd1 vccd1 vccd1 _12473_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10490_ _12495_/Q _12494_/Q _09135_/B vssd1 vssd1 vccd1 vccd1 _10490_/X sky130_fd_sc_hd__a21bo_1
XFILLER_136_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09149_ _12594_/Q vssd1 vssd1 vccd1 vccd1 _09175_/B sky130_fd_sc_hd__inv_2
XFILLER_136_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12160_ _10784_/X _11142_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _12160_/X sky130_fd_sc_hd__mux2_2
XFILLER_146_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11111_ _11111_/A vssd1 vssd1 vccd1 vccd1 _11111_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12091_ _12448_/Q _12090_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _12091_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11042_ _06392_/X _10691_/A _11032_/X _11041_/X _11034_/X vssd1 vssd1 vccd1 vccd1
+ _11042_/X sky130_fd_sc_hd__a32o_1
XFILLER_104_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12993_ _12993_/CLK _12993_/D vssd1 vssd1 vccd1 vccd1 _12993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11944_ _09720_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11944_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11875_ _10278_/X _12816_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11875_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10826_ _12516_/Q _12328_/Q _10824_/Y _10825_/Y vssd1 vssd1 vccd1 vccd1 _10827_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_60_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10757_ _12763_/Q _12762_/Q vssd1 vssd1 vccd1 vccd1 _10757_/Y sky130_fd_sc_hd__nor2_2
XFILLER_13_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10688_ _06410_/X _11034_/A _10686_/X _11045_/A vssd1 vssd1 vccd1 vccd1 _10688_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_187_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12427_ _12471_/CLK _12427_/D vssd1 vssd1 vccd1 vccd1 _12427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12358_ _13257_/CLK _12358_/D vssd1 vssd1 vccd1 vccd1 _12358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11309_ vssd1 vssd1 vccd1 vccd1 _11309_/HI _11309_/LO sky130_fd_sc_hd__conb_1
XFILLER_114_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12289_ _12296_/CLK _12289_/D vssd1 vssd1 vccd1 vccd1 _12289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06850_ _06848_/X _06849_/X _06848_/X _06849_/X vssd1 vssd1 vccd1 vccd1 _06850_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06781_ _12004_/X _06760_/X _12004_/X _06760_/X vssd1 vssd1 vccd1 vccd1 _06783_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08520_ _08519_/X _12248_/X _08514_/X _12761_/Q vssd1 vssd1 vccd1 vccd1 _12761_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08451_ _13073_/Q _07809_/Y _13055_/Q _10352_/A vssd1 vssd1 vccd1 vccd1 _08451_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07402_ _07408_/A vssd1 vssd1 vccd1 vccd1 _07402_/X sky130_fd_sc_hd__clkbuf_1
X_08382_ _12794_/Q _08374_/X _08005_/X _08375_/X vssd1 vssd1 vccd1 vccd1 _12794_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07333_ _07345_/A vssd1 vssd1 vccd1 vccd1 _07333_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_118_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 _12718_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07264_ _07264_/A vssd1 vssd1 vccd1 vccd1 _07264_/X sky130_fd_sc_hd__buf_2
XFILLER_191_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09003_ _09019_/B vssd1 vssd1 vccd1 vccd1 _09008_/B sky130_fd_sc_hd__clkbuf_2
X_06215_ _13280_/Q vssd1 vssd1 vccd1 vccd1 _06215_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07195_ _11964_/S vssd1 vssd1 vccd1 vccd1 _09982_/B sky130_fd_sc_hd__buf_2
XFILLER_191_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06146_ _12742_/Q _12710_/Q _12741_/Q _12709_/Q vssd1 vssd1 vccd1 vccd1 _06146_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06077_ _12730_/Q _12698_/Q _06076_/X vssd1 vssd1 vccd1 vccd1 _06077_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_132_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09905_ _09903_/Y _09897_/X _06332_/A _09892_/X _09904_/X vssd1 vssd1 vccd1 vccd1
+ _09905_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09836_ _13231_/Q vssd1 vssd1 vccd1 vccd1 _09836_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09767_ _09764_/Y _09766_/A _09769_/B _09766_/Y _09492_/A vssd1 vssd1 vccd1 vccd1
+ _09768_/B sky130_fd_sc_hd__o221a_1
XFILLER_86_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06979_ _06841_/A _06971_/B _06977_/Y _06630_/X _09550_/B vssd1 vssd1 vccd1 vccd1
+ _06980_/A sky130_fd_sc_hd__o32a_1
XFILLER_67_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08729_/A sky130_fd_sc_hd__clkbuf_2
XPHY_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09698_ _09698_/A vssd1 vssd1 vccd1 vccd1 _09698_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _08653_/A vssd1 vssd1 vccd1 vccd1 _08649_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_199_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11660_ _11659_/X _10522_/Y _11704_/S vssd1 vssd1 vccd1 vccd1 _12372_/D sky130_fd_sc_hd__mux2_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10611_ _10611_/A _10611_/B vssd1 vssd1 vccd1 vccd1 _10612_/A sky130_fd_sc_hd__or2_1
XPHY_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ _10438_/X _09244_/A _11592_/S vssd1 vssd1 vccd1 vccd1 _11591_/X sky130_fd_sc_hd__mux2_1
XPHY_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10542_ _09329_/A _09329_/B _10541_/Y vssd1 vssd1 vccd1 vccd1 _10542_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _13264_/CLK _13261_/D _06319_/X vssd1 vssd1 vccd1 vccd1 _13261_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10473_ _08164_/Y _10468_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _10474_/C sky130_fd_sc_hd__o21a_1
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ _12211_/X _12626_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12212_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ _13237_/CLK _13192_/D _06843_/X vssd1 vssd1 vccd1 vccd1 _13192_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_159_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12143_ _12142_/X _12438_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12143_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12074_ _12446_/Q _12073_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _12074_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11025_ _11024_/A _11024_/B _12321_/D vssd1 vssd1 vccd1 vccd1 _12361_/D sky130_fd_sc_hd__a21oi_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12976_ _12976_/CLK _12976_/D vssd1 vssd1 vccd1 vccd1 _12976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11927_ _09480_/X _12788_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11927_/X sky130_fd_sc_hd__mux2_2
XPHY_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11858_ _10069_/Y _12314_/Q _12312_/Q vssd1 vssd1 vccd1 vccd1 _11858_/X sky130_fd_sc_hd__mux2_2
XFILLER_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10809_ _12512_/Q _12324_/Q _10806_/Y _10804_/Y vssd1 vssd1 vccd1 vccd1 _10809_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_11789_ _12130_/X _11788_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11789_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07951_ _07951_/A vssd1 vssd1 vccd1 vccd1 _07962_/S sky130_fd_sc_hd__buf_2
XFILLER_141_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06902_ _06900_/X _06901_/X _06900_/X _06901_/X vssd1 vssd1 vccd1 vccd1 _06902_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07882_ _12840_/Q _07888_/A _07881_/Y vssd1 vssd1 vccd1 vccd1 _10324_/A sky130_fd_sc_hd__o21ai_4
XFILLER_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06833_ _06831_/X _06832_/X _06831_/X _06832_/X vssd1 vssd1 vccd1 vccd1 _06840_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_09621_ _09620_/A _09620_/B _09643_/A vssd1 vssd1 vccd1 vccd1 _09621_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09552_ _09552_/A _09552_/B _09552_/C vssd1 vssd1 vccd1 vccd1 _09566_/A sky130_fd_sc_hd__nor3_4
X_06764_ _06630_/X _06754_/X _06762_/X _06646_/X _06763_/Y vssd1 vssd1 vccd1 vccd1
+ _06765_/A sky130_fd_sc_hd__a32o_1
XFILLER_110_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08503_ _08503_/A vssd1 vssd1 vccd1 vccd1 _08503_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09483_ _09482_/A _09482_/B _09482_/C vssd1 vssd1 vccd1 vccd1 _09483_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_93_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06695_ _12756_/Q vssd1 vssd1 vccd1 vccd1 _11034_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08434_ _12774_/Q _08417_/A _07564_/X _08418_/A vssd1 vssd1 vccd1 vccd1 _12774_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08365_ _12801_/Q _08358_/X _07983_/X _08360_/X vssd1 vssd1 vccd1 vccd1 _12801_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07316_ _09071_/C _09072_/A _09071_/D vssd1 vssd1 vccd1 vccd1 _09042_/B sky130_fd_sc_hd__or3b_1
XFILLER_149_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08296_ _08296_/A vssd1 vssd1 vccd1 vccd1 _08296_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07247_ _07251_/A vssd1 vssd1 vccd1 vccd1 _07247_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_165_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07178_ _11522_/X _07176_/X _13121_/Q _07177_/X vssd1 vssd1 vccd1 vccd1 _13121_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06129_ _06129_/A vssd1 vssd1 vccd1 vccd1 _06130_/C sky130_fd_sc_hd__inv_2
XFILLER_105_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_86_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _12769_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09819_ _09886_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09819_/X sky130_fd_sc_hd__or2_1
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12830_ _12169_/X _12830_/D _08291_/X vssd1 vssd1 vccd1 vccd1 _12830_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12761_ _12986_/CLK _12761_/D _08518_/X vssd1 vssd1 vccd1 vccd1 _12761_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11712_ _11711_/X _10638_/Y _11774_/S vssd1 vssd1 vccd1 vccd1 _12420_/D sky130_fd_sc_hd__mux2_1
XPHY_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12725_/CLK _12692_/D _08723_/X vssd1 vssd1 vccd1 vccd1 _12692_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_199_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11643_ _10513_/X _12928_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11643_/X sky130_fd_sc_hd__mux2_1
XPHY_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11574_ _12831_/Q _10794_/C _11578_/S vssd1 vssd1 vccd1 vccd1 _11574_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput17 io_in[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_1
XFILLER_195_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 io_in[34] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
XFILLER_183_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10525_ _10525_/A _10586_/A _10585_/A _10525_/D vssd1 vssd1 vccd1 vccd1 _10526_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_11_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput39 la_data_in[0] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_4
XPHY_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13244_ _13244_/CLK _13244_/D _06391_/X vssd1 vssd1 vccd1 vccd1 _13244_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_170_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10456_ _10460_/B vssd1 vssd1 vccd1 vccd1 _10463_/C sky130_fd_sc_hd__inv_2
X_13175_ _13183_/CLK _13175_/D _06985_/X vssd1 vssd1 vccd1 vccd1 _13175_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10387_ _10387_/A _10388_/B _10387_/C vssd1 vssd1 vccd1 vccd1 _10387_/Y sky130_fd_sc_hd__nor3_1
XFILLER_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12126_ _12437_/Q _10675_/Y _12139_/S vssd1 vssd1 vccd1 vccd1 _12126_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12057_ _12056_/X _12439_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__mux2_1
Xrepeater607 _11634_/S vssd1 vssd1 vccd1 vccd1 _12307_/D sky130_fd_sc_hd__clkbuf_8
Xrepeater618 _11487_/S vssd1 vssd1 vccd1 vccd1 _11492_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater629 _11546_/S vssd1 vssd1 vccd1 vccd1 _11543_/S sky130_fd_sc_hd__buf_6
X_11008_ _12355_/Q _11004_/Y _11010_/A vssd1 vssd1 vccd1 vccd1 _12355_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12959_ _12976_/CLK _12959_/D vssd1 vssd1 vccd1 vccd1 _12959_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06480_ _06841_/A vssd1 vssd1 vccd1 vccd1 _06480_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_179_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08150_ _13128_/Q _10444_/B _13142_/Q _10480_/A vssd1 vssd1 vccd1 vccd1 _08150_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07101_ _07101_/A _07101_/B _07101_/C _07101_/D vssd1 vssd1 vccd1 vccd1 _07102_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08081_ _08085_/A vssd1 vssd1 vccd1 vccd1 _08081_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07032_ _07046_/A vssd1 vssd1 vccd1 vccd1 _07032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ _07508_/Y _07512_/Y _09284_/C _12572_/Q vssd1 vssd1 vccd1 vccd1 _09279_/D
+ sky130_fd_sc_hd__a31o_1
X_07934_ _07945_/A vssd1 vssd1 vccd1 vccd1 _07934_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07865_ _13020_/Q _10346_/A _07820_/Y _07821_/X vssd1 vssd1 vccd1 vccd1 _07866_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09604_ _09604_/A _09604_/B _09604_/C vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__nor3_4
X_06816_ _12019_/X _12018_/X _06815_/X vssd1 vssd1 vccd1 vccd1 _06816_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07796_ _12897_/Q vssd1 vssd1 vccd1 vccd1 _10328_/A sky130_fd_sc_hd__inv_2
XFILLER_113_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06747_ _06750_/A vssd1 vssd1 vccd1 vccd1 _06747_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09535_ _13153_/Q vssd1 vssd1 vccd1 vccd1 _09535_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_133_wb_clk_i _12726_/CLK vssd1 vssd1 vccd1 vccd1 _12688_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ _12604_/Q _07518_/A _13008_/Q _09442_/A vssd1 vssd1 vccd1 vccd1 _09466_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06678_ _06665_/X _06669_/X _06671_/Y vssd1 vssd1 vccd1 vccd1 _06678_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08417_ _08417_/A vssd1 vssd1 vccd1 vccd1 _08417_/X sky130_fd_sc_hd__clkbuf_2
X_09397_ _09362_/Y _12398_/D _12459_/Q _10521_/A _09396_/X vssd1 vssd1 vccd1 vccd1
+ _09402_/C sky130_fd_sc_hd__o221a_1
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08348_ _08352_/A vssd1 vssd1 vccd1 vccd1 _08348_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_184_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08279_ _08337_/A vssd1 vssd1 vccd1 vccd1 _08353_/S sky130_fd_sc_hd__clkbuf_4
X_10310_ _13270_/Q vssd1 vssd1 vccd1 vccd1 _10310_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11290_ vssd1 vssd1 vccd1 vccd1 _11290_/HI _11290_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10241_ _10237_/Y _10163_/X _10238_/Y _10165_/X _10240_/X vssd1 vssd1 vccd1 vccd1
+ _10241_/X sky130_fd_sc_hd__o221a_1
XFILLER_98_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10172_ _09909_/Y _10134_/X _10159_/X _10171_/X vssd1 vssd1 vccd1 vccd1 _10172_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_120_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput490 _11240_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12813_ _12169_/X _12813_/D _08332_/X vssd1 vssd1 vccd1 vccd1 _12813_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12744_ _12747_/CLK _12744_/D _08589_/X vssd1 vssd1 vccd1 vccd1 _12744_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_76_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12679_/CLK _12675_/D _08776_/X vssd1 vssd1 vccd1 vccd1 _12675_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _10496_/X _12993_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11626_/X sky130_fd_sc_hd__mux2_1
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11557_ _12814_/Q _09243_/C _11558_/S vssd1 vssd1 vccd1 vccd1 _11557_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10508_ _12582_/Q _07756_/B _07757_/B vssd1 vssd1 vccd1 vccd1 _10508_/X sky130_fd_sc_hd__a21bo_1
X_11488_ _10334_/Y _09184_/B _11492_/S vssd1 vssd1 vccd1 vccd1 _11488_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13227_ _13227_/CLK _13227_/D _06506_/X vssd1 vssd1 vccd1 vccd1 _13227_/Q sky130_fd_sc_hd__dfrtp_1
X_10439_ _10439_/A _10439_/B _10439_/C vssd1 vssd1 vccd1 vccd1 _10444_/C sky130_fd_sc_hd__or3_4
XFILLER_83_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13158_ _13158_/CLK _13158_/D _07052_/X vssd1 vssd1 vccd1 vccd1 _13158_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12109_ _12432_/Q _10669_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12109_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13089_ _12167_/X _13089_/D _07262_/X vssd1 vssd1 vccd1 vccd1 _13089_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07650_ _07661_/A _07650_/B _07658_/A _07650_/D vssd1 vssd1 vccd1 vccd1 _07651_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06601_ _06650_/A vssd1 vssd1 vccd1 vccd1 _06601_/X sky130_fd_sc_hd__clkbuf_1
X_07581_ _12981_/Q _07574_/X _07562_/A _07575_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _12981_/D sky130_fd_sc_hd__o221a_1
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09320_ _12369_/Q vssd1 vssd1 vccd1 vccd1 _09332_/A sky130_fd_sc_hd__inv_2
X_06532_ _06580_/A vssd1 vssd1 vccd1 vccd1 _06532_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ _09251_/A vssd1 vssd1 vccd1 vccd1 _09251_/X sky130_fd_sc_hd__clkbuf_2
X_06463_ _06444_/A _06444_/B _06444_/Y vssd1 vssd1 vccd1 vccd1 _06463_/Y sky130_fd_sc_hd__a21oi_1
X_08202_ _13092_/Q vssd1 vssd1 vccd1 vccd1 _08202_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09182_ _09243_/A _10528_/C _09244_/A _09244_/B vssd1 vssd1 vccd1 vccd1 _09183_/D
+ sky130_fd_sc_hd__or4_4
X_06394_ _06416_/A vssd1 vssd1 vccd1 vccd1 _06412_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08133_ _12826_/Q vssd1 vssd1 vccd1 vccd1 _10467_/B sky130_fd_sc_hd__inv_2
XFILLER_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08064_ _10035_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08067_/A sky130_fd_sc_hd__or2_1
XFILLER_190_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07015_ _06886_/X _12186_/X _06887_/X _13170_/Q vssd1 vssd1 vccd1 vccd1 _13170_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_175_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput207 la_oenb[20] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__buf_1
Xinput218 la_oenb[30] vssd1 vssd1 vccd1 vccd1 input218/X sky130_fd_sc_hd__buf_1
Xinput229 la_oenb[40] vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_hd__buf_1
X_08966_ _08969_/A vssd1 vssd1 vccd1 vccd1 _08966_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07917_ _07917_/A vssd1 vssd1 vccd1 vccd1 _07917_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08897_ _08897_/A vssd1 vssd1 vccd1 vccd1 _08897_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07848_ _13029_/Q _10373_/A _13024_/Q _10357_/A vssd1 vssd1 vccd1 vccd1 _07848_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07779_ _07781_/A vssd1 vssd1 vccd1 vccd1 _07780_/A sky130_fd_sc_hd__inv_2
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09518_ _09502_/X _09505_/Y _09516_/Y _09492_/A _09517_/Y vssd1 vssd1 vccd1 vccd1
+ _09518_/X sky130_fd_sc_hd__o311a_1
XFILLER_140_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10790_ _10790_/A vssd1 vssd1 vccd1 vccd1 _10790_/Y sky130_fd_sc_hd__inv_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _12979_/Q _09436_/X _12927_/Q _09438_/X _09448_/X vssd1 vssd1 vccd1 vccd1
+ _09449_/X sky130_fd_sc_hd__a221o_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _12978_/CLK _12460_/D vssd1 vssd1 vccd1 vccd1 _12460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11411_ _11410_/X _12443_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _11411_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12391_ _12413_/CLK _12391_/D vssd1 vssd1 vccd1 vccd1 _12413_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_153_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11342_ vssd1 vssd1 vccd1 vccd1 _11342_/HI _11342_/LO sky130_fd_sc_hd__conb_1
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12620_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11273_ vssd1 vssd1 vccd1 vccd1 _11273_/HI _11273_/LO sky130_fd_sc_hd__conb_1
XFILLER_125_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13012_ _12164_/X _13012_/D _07485_/X vssd1 vssd1 vccd1 vccd1 _13012_/Q sky130_fd_sc_hd__dfrtp_1
X_10224_ _10219_/Y _10163_/X _10220_/Y _10165_/X _10223_/X vssd1 vssd1 vccd1 vccd1
+ _10224_/X sky130_fd_sc_hd__o221a_1
XFILLER_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10155_ _07869_/Y _10151_/X _10154_/X vssd1 vssd1 vccd1 vccd1 _10155_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_94_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10086_ _10792_/D _10035_/A _10084_/Y _10085_/Y _10140_/A vssd1 vssd1 vccd1 vccd1
+ _10086_/X sky130_fd_sc_hd__o32a_1
XFILLER_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10988_ _11000_/C vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12727_ _12737_/CLK _12727_/D _08634_/X vssd1 vssd1 vccd1 vccd1 _12727_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ _13264_/CLK _12658_/D _08826_/X vssd1 vssd1 vccd1 vccd1 _12658_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11609_ _10485_/X _10793_/B _11610_/S vssd1 vssd1 vccd1 vccd1 _11609_/X sky130_fd_sc_hd__mux2_1
X_12589_ _12937_/CLK _12589_/D vssd1 vssd1 vccd1 vccd1 _12589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08820_ _08814_/X _08817_/X _06316_/X _12661_/Q _08811_/X vssd1 vssd1 vccd1 vccd1
+ _12661_/D sky130_fd_sc_hd__a32o_1
XFILLER_98_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08751_ _08839_/A vssd1 vssd1 vccd1 vccd1 _08769_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07702_ _07702_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07702_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08682_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08682_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07633_ _12951_/Q _12950_/Q _07658_/A _07650_/B vssd1 vssd1 vccd1 vccd1 _07660_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07564_ _09226_/A vssd1 vssd1 vccd1 vccd1 _07564_/X sky130_fd_sc_hd__buf_4
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09303_ _10655_/B vssd1 vssd1 vccd1 vccd1 _11818_/S sky130_fd_sc_hd__inv_16
X_06515_ _06509_/Y _06510_/Y _06549_/A _06514_/X vssd1 vssd1 vccd1 vccd1 _06520_/A
+ sky130_fd_sc_hd__a31o_1
X_07495_ _07775_/A vssd1 vssd1 vccd1 vccd1 _07609_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _12466_/Q _09231_/X _07545_/X _09233_/X vssd1 vssd1 vccd1 vccd1 _12466_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06446_ _10714_/B _06446_/B vssd1 vssd1 vccd1 vccd1 _10711_/A sky130_fd_sc_hd__or2_2
XFILLER_107_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09165_ _11628_/X _09163_/X _12503_/Q _09164_/X vssd1 vssd1 vccd1 vccd1 _12503_/D
+ sky130_fd_sc_hd__a22o_1
X_06377_ _06361_/X _12224_/X _06375_/X _06376_/X vssd1 vssd1 vccd1 vccd1 _13249_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_194_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08116_ _13121_/Q vssd1 vssd1 vccd1 vccd1 _08116_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09096_ _12538_/Q _09089_/X _10794_/B _09092_/X vssd1 vssd1 vccd1 vccd1 _12538_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08047_ _08051_/A vssd1 vssd1 vccd1 vccd1 _08047_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_190_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09998_ _08777_/Y _09993_/X _06236_/Y _09972_/X _09991_/X vssd1 vssd1 vccd1 vccd1
+ _09998_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_77_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08949_ _09312_/A _08949_/B vssd1 vssd1 vccd1 vccd1 _12140_/S sky130_fd_sc_hd__or2_4
XFILLER_29_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11960_ _09267_/X _09266_/Y _12549_/Q vssd1 vssd1 vccd1 vccd1 _12549_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10911_ _12529_/Q vssd1 vssd1 vccd1 vccd1 _10911_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11891_ _08926_/A _10633_/X _12321_/Q vssd1 vssd1 vccd1 vccd1 _11891_/X sky130_fd_sc_hd__mux2_1
X_10842_ _12331_/Q vssd1 vssd1 vccd1 vccd1 _10843_/B sky130_fd_sc_hd__inv_2
XFILLER_60_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10773_ _10773_/A vssd1 vssd1 vccd1 vccd1 _10773_/X sky130_fd_sc_hd__buf_2
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12512_ _12517_/CLK _12512_/D vssd1 vssd1 vccd1 vccd1 _12512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12443_ _12489_/CLK _12443_/D vssd1 vssd1 vccd1 vccd1 _12443_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12374_ _12376_/CLK _12374_/D vssd1 vssd1 vccd1 vccd1 _12396_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_176_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11325_ vssd1 vssd1 vccd1 vccd1 _11325_/HI _11325_/LO sky130_fd_sc_hd__conb_1
XFILLER_158_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11256_ vssd1 vssd1 vccd1 vccd1 _11256_/HI _11256_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10207_ _10227_/A _11980_/X vssd1 vssd1 vccd1 vccd1 _10207_/Y sky130_fd_sc_hd__nor2b_4
X_11187_ vssd1 vssd1 vccd1 vccd1 _11187_/HI _11187_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10138_ _10135_/Y _10000_/A _10136_/Y _10137_/X vssd1 vssd1 vccd1 vccd1 _10138_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10069_ _10150_/A _11973_/X vssd1 vssd1 vccd1 vccd1 _10069_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_169_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06300_ _06300_/A vssd1 vssd1 vccd1 vccd1 _06300_/Y sky130_fd_sc_hd__clkinv_4
X_07280_ _07280_/A vssd1 vssd1 vccd1 vccd1 _07280_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06231_ _13277_/Q vssd1 vssd1 vccd1 vccd1 _06231_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06162_ _06162_/A vssd1 vssd1 vccd1 vccd1 _06217_/A sky130_fd_sc_hd__buf_2
XFILLER_117_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06093_ _12726_/Q _12694_/Q _12725_/Q _12693_/Q vssd1 vssd1 vccd1 vccd1 _06093_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09921_ _12664_/Q vssd1 vssd1 vccd1 vccd1 _09921_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09852_ _09803_/X _09851_/B _09849_/Y _09881_/A _09851_/X vssd1 vssd1 vccd1 vccd1
+ _09854_/B sky130_fd_sc_hd__o311a_1
XFILLER_86_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08803_ _08807_/A vssd1 vssd1 vccd1 vccd1 _08803_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09783_ _09782_/A _09782_/B _09782_/Y vssd1 vssd1 vccd1 vccd1 _09802_/A sky130_fd_sc_hd__a21o_1
XFILLER_26_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06995_ _06995_/A _06995_/B vssd1 vssd1 vccd1 vccd1 _06995_/X sky130_fd_sc_hd__or2_1
XFILLER_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08734_ _08747_/A vssd1 vssd1 vccd1 vccd1 _08734_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _08669_/A vssd1 vssd1 vccd1 vccd1 _08665_/X sky130_fd_sc_hd__clkbuf_1
XPHY_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _09009_/A vssd1 vssd1 vccd1 vccd1 _07616_/X sky130_fd_sc_hd__clkbuf_4
XPHY_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _08606_/A vssd1 vssd1 vccd1 vccd1 _08596_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07547_ _07547_/A vssd1 vssd1 vccd1 vccd1 _09441_/A sky130_fd_sc_hd__inv_2
XFILLER_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07478_ _07933_/A vssd1 vssd1 vccd1 vccd1 _07489_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09217_ _12474_/Q _09215_/X _07558_/X _09216_/X vssd1 vssd1 vccd1 vccd1 _12474_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06429_ _12131_/X vssd1 vssd1 vccd1 vccd1 _06430_/A sky130_fd_sc_hd__inv_2
XFILLER_167_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09148_ _12965_/Q vssd1 vssd1 vccd1 vccd1 _09150_/A sky130_fd_sc_hd__inv_2
XFILLER_147_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09079_ _09079_/A vssd1 vssd1 vccd1 vccd1 _09079_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11110_ _11110_/A vssd1 vssd1 vccd1 vccd1 _11110_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12090_ _12448_/Q _10684_/X _12090_/S vssd1 vssd1 vccd1 vccd1 _12090_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11041_ _11041_/A vssd1 vssd1 vccd1 vccd1 _11041_/X sky130_fd_sc_hd__buf_2
XFILLER_118_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12992_ _12992_/CLK _12992_/D vssd1 vssd1 vccd1 vccd1 _12992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11943_ _09700_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11943_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11874_ _10261_/X _12815_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11874_/X sky130_fd_sc_hd__mux2_1
X_10825_ _12328_/Q vssd1 vssd1 vccd1 vccd1 _10825_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10756_ _10755_/X _10750_/X _06371_/X _10751_/X _10752_/X vssd1 vssd1 vccd1 vccd1
+ _10756_/X sky130_fd_sc_hd__a221o_1
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ _10687_/A vssd1 vssd1 vccd1 vccd1 _11045_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_199_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12426_ _12426_/CLK _12426_/D vssd1 vssd1 vccd1 vccd1 _12426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12357_ _12357_/CLK _12357_/D vssd1 vssd1 vccd1 vccd1 _12357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ vssd1 vssd1 vccd1 vccd1 _11308_/HI _11308_/LO sky130_fd_sc_hd__conb_1
XFILLER_113_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12288_ _12296_/CLK _12288_/D vssd1 vssd1 vccd1 vccd1 _12288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11239_ vssd1 vssd1 vccd1 vccd1 _11239_/HI _11239_/LO sky130_fd_sc_hd__conb_1
XFILLER_68_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06780_ _06806_/A vssd1 vssd1 vccd1 vccd1 _06780_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08450_ _13052_/Q vssd1 vssd1 vccd1 vccd1 _08450_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07401_ _11418_/X _07368_/A _13042_/Q _07369_/A vssd1 vssd1 vccd1 vccd1 _13042_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08381_ _08385_/A vssd1 vssd1 vccd1 vccd1 _08381_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07332_ _07362_/A vssd1 vssd1 vccd1 vccd1 _07345_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07263_ _07263_/A vssd1 vssd1 vccd1 vccd1 _07263_/X sky130_fd_sc_hd__buf_2
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09002_ _09002_/A _12595_/Q vssd1 vssd1 vccd1 vccd1 _12593_/D sky130_fd_sc_hd__or2_1
X_06214_ _06214_/A vssd1 vssd1 vccd1 vccd1 _06214_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07194_ _07206_/A vssd1 vssd1 vccd1 vccd1 _07194_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06145_ _06144_/A _06070_/X _06134_/Y _06197_/A _06144_/X vssd1 vssd1 vccd1 vccd1
+ _06145_/X sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_158_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12529_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_191_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06076_ _12730_/Q _12698_/Q _12729_/Q _12697_/Q vssd1 vssd1 vccd1 vccd1 _06076_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09904_ _12881_/Q _09910_/B vssd1 vssd1 vccd1 vccd1 _09904_/X sky130_fd_sc_hd__or2_1
XFILLER_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09835_ _13230_/Q _13229_/Q _06483_/Y _06488_/Y vssd1 vssd1 vccd1 vccd1 _09837_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_59_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09766_ _09766_/A vssd1 vssd1 vccd1 vccd1 _09766_/Y sky130_fd_sc_hd__inv_2
X_06978_ _13177_/Q vssd1 vssd1 vccd1 vccd1 _09550_/B sky130_fd_sc_hd__inv_2
XPHY_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08717_ _11829_/X _08715_/X _12695_/Q _08716_/X vssd1 vssd1 vccd1 vccd1 _12695_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _09671_/A _09671_/B _09677_/X vssd1 vssd1 vccd1 vccd1 _09698_/A sky130_fd_sc_hd__o21ai_1
XPHY_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08648_ _11931_/X _08639_/X _12722_/Q _08640_/X vssd1 vssd1 vccd1 vccd1 _12722_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _11958_/X _08575_/X _12749_/Q _08578_/X vssd1 vssd1 vccd1 vccd1 _12749_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10610_ _12415_/D _10610_/B _12413_/D _12414_/D vssd1 vssd1 vccd1 vccd1 _11406_/S
+ sky130_fd_sc_hd__or4_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11590_ _10436_/Y _09244_/B _11592_/S vssd1 vssd1 vccd1 vccd1 _11590_/X sky130_fd_sc_hd__mux2_1
XPHY_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10541_ _10541_/A vssd1 vssd1 vccd1 vccd1 _10541_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ _13260_/CLK _13260_/D _06325_/X vssd1 vssd1 vccd1 vccd1 _13260_/Q sky130_fd_sc_hd__dfrtp_1
X_10472_ _12829_/Q _12828_/Q _10472_/C vssd1 vssd1 vccd1 vccd1 _10475_/B sky130_fd_sc_hd__and3_1
X_12211_ _06332_/Y _13151_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12211_/X sky130_fd_sc_hd__mux2_1
X_13191_ _13193_/CLK _13191_/D _06859_/X vssd1 vssd1 vccd1 vccd1 _13191_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12142_ _12141_/X _12438_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12142_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12073_ _12446_/Q _10682_/X _12090_/S vssd1 vssd1 vccd1 vccd1 _12073_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11024_ _11024_/A _11024_/B vssd1 vssd1 vccd1 vccd1 _12321_/D sky130_fd_sc_hd__nor2_1
XFILLER_1_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12975_ _12975_/CLK _12975_/D vssd1 vssd1 vccd1 vccd1 _12975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _12844_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_11926_ _10311_/Y _12803_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _11926_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11857_ _10072_/Y _12805_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11857_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10808_ _10806_/A _10807_/A _10806_/Y _10807_/Y vssd1 vssd1 vccd1 vccd1 _12324_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11788_ _09244_/A _11787_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11788_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10739_ _12131_/X vssd1 vssd1 vccd1 vccd1 _10739_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12409_ _12458_/CLK _12409_/D vssd1 vssd1 vccd1 vccd1 _12409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07950_ _07961_/A vssd1 vssd1 vccd1 vccd1 _07950_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06901_ _12024_/X _12020_/X _12024_/X _12020_/X vssd1 vssd1 vccd1 vccd1 _06901_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07881_ _12842_/Q vssd1 vssd1 vccd1 vccd1 _07881_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09620_ _09620_/A _09620_/B vssd1 vssd1 vccd1 vccd1 _09643_/A sky130_fd_sc_hd__or2_2
X_06832_ _06813_/A _06813_/B _06813_/X vssd1 vssd1 vccd1 vccd1 _06832_/X sky130_fd_sc_hd__a21bo_1
XFILLER_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09551_ _09550_/A _09550_/B _09550_/Y vssd1 vssd1 vccd1 vccd1 _09552_/C sky130_fd_sc_hd__a21o_1
X_06763_ _13202_/Q vssd1 vssd1 vccd1 vccd1 _06763_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08502_ _06403_/X _12262_/X _08499_/X _12768_/Q vssd1 vssd1 vccd1 vccd1 _12768_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06694_ _06694_/A _06694_/B vssd1 vssd1 vccd1 vccd1 _06694_/X sky130_fd_sc_hd__or2_1
X_09482_ _09482_/A _09482_/B _09482_/C vssd1 vssd1 vccd1 vccd1 _09487_/A sky130_fd_sc_hd__or3_1
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08433_ _08433_/A vssd1 vssd1 vccd1 vccd1 _08433_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08364_ _08370_/A vssd1 vssd1 vccd1 vccd1 _08364_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07315_ _07330_/A vssd1 vssd1 vccd1 vccd1 _07315_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08295_ _12829_/Q _11604_/X _08307_/S vssd1 vssd1 vccd1 vccd1 _12829_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07246_ _11561_/X _07233_/X _13096_/Q _07234_/X vssd1 vssd1 vccd1 vccd1 _13096_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07177_ _07177_/A vssd1 vssd1 vccd1 vccd1 _07177_/X sky130_fd_sc_hd__buf_2
XFILLER_173_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06128_ _06174_/A _06175_/B _06174_/A _06175_/A _06176_/A vssd1 vssd1 vccd1 vccd1
+ _06129_/A sky130_fd_sc_hd__o221a_1
XFILLER_133_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06059_ _12735_/Q _12703_/Q _12735_/Q _12703_/Q vssd1 vssd1 vccd1 vccd1 _06259_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09818_ _09823_/B _09817_/Y _09815_/A _09817_/A _09492_/A vssd1 vssd1 vccd1 vccd1
+ _09819_/B sky130_fd_sc_hd__o221a_1
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_wb_clk_i _12328_/CLK vssd1 vssd1 vccd1 vccd1 _12779_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09749_ _09709_/Y _09711_/Y _09729_/Y vssd1 vssd1 vccd1 vccd1 _09749_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12760_ _12986_/CLK _12760_/D _08522_/X vssd1 vssd1 vccd1 vccd1 _12760_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_199_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11711_ _10638_/Y _10639_/Y _11818_/S vssd1 vssd1 vccd1 vccd1 _11711_/X sky130_fd_sc_hd__mux2_1
XPHY_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12725_/CLK _12691_/D _08725_/X vssd1 vssd1 vccd1 vccd1 _12691_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _10512_/X _12927_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11642_/X sky130_fd_sc_hd__mux2_1
XPHY_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11573_ _12830_/Q _10794_/D _11578_/S vssd1 vssd1 vccd1 vccd1 _11573_/X sky130_fd_sc_hd__mux2_1
XPHY_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 io_in[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_1
XPHY_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput29 io_in[35] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
XFILLER_196_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10524_ _10603_/A _12410_/D _10599_/A _12408_/D vssd1 vssd1 vccd1 vccd1 _10525_/D
+ sky130_fd_sc_hd__or4_4
XPHY_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13243_ _13243_/CLK _13243_/D _06395_/X vssd1 vssd1 vccd1 vccd1 _13243_/Q sky130_fd_sc_hd__dfrtp_2
X_10455_ _10455_/A _10455_/B _10455_/C _10455_/D vssd1 vssd1 vccd1 vccd1 _10460_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_184_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13174_ _13177_/CLK _13174_/D _06994_/X vssd1 vssd1 vccd1 vccd1 _13174_/Q sky130_fd_sc_hd__dfrtp_1
X_10386_ _07868_/Y _10381_/A _07824_/Y vssd1 vssd1 vccd1 vccd1 _10387_/C sky130_fd_sc_hd__o21a_1
X_12125_ _12124_/X _12434_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12125_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12056_ _12439_/Q _10677_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _12056_/X sky130_fd_sc_hd__mux2_1
Xrepeater608 _11348_/X vssd1 vssd1 vccd1 vccd1 _12282_/S0 sky130_fd_sc_hd__buf_12
Xrepeater619 _11469_/S vssd1 vssd1 vccd1 vccd1 _11481_/S sky130_fd_sc_hd__buf_6
X_11007_ _11014_/A _11014_/B _11014_/D vssd1 vssd1 vccd1 vccd1 _11010_/A sky130_fd_sc_hd__or3_4
XFILLER_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12958_ _12961_/CLK _12958_/D vssd1 vssd1 vccd1 vccd1 _12958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11909_ _11908_/X _12142_/S _11909_/S vssd1 vssd1 vccd1 vccd1 _11909_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12889_ _12890_/CLK _12889_/D _07985_/X vssd1 vssd1 vccd1 vccd1 _12889_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07100_ _07100_/A _07100_/B vssd1 vssd1 vccd1 vccd1 _07102_/C sky130_fd_sc_hd__nand2_1
XFILLER_201_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08080_ _12855_/Q _08066_/X _07993_/X _08068_/X vssd1 vssd1 vccd1 vccd1 _12855_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07031_ _06663_/X _07030_/X _06415_/B _13164_/Q vssd1 vssd1 vccd1 vccd1 _13164_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_162_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08982_ _12299_/Q vssd1 vssd1 vccd1 vccd1 _09279_/A sky130_fd_sc_hd__inv_2
XFILLER_115_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07933_ _07933_/A vssd1 vssd1 vccd1 vccd1 _07945_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07864_ _13027_/Q _10367_/B _13020_/Q _10346_/A vssd1 vssd1 vccd1 vccd1 _07866_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_29_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09603_ _13188_/Q _09602_/B _09614_/A vssd1 vssd1 vccd1 vccd1 _09604_/C sky130_fd_sc_hd__o21ai_2
X_06815_ _12010_/X _06815_/B vssd1 vssd1 vccd1 vccd1 _06815_/X sky130_fd_sc_hd__or2_1
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07795_ _13011_/Q vssd1 vssd1 vccd1 vccd1 _07795_/Y sky130_fd_sc_hd__inv_2
X_09534_ _09530_/X _09531_/Y _09533_/X vssd1 vssd1 vccd1 vccd1 _09534_/Y sky130_fd_sc_hd__o21ai_1
X_06746_ _06658_/X _06739_/Y _06608_/X _06745_/X vssd1 vssd1 vccd1 vccd1 _13204_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09465_ _12984_/Q _09436_/X _13007_/Q _09442_/X _09464_/X vssd1 vssd1 vccd1 vccd1
+ _09465_/X sky130_fd_sc_hd__a221o_1
XPHY_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06677_ _13211_/Q vssd1 vssd1 vccd1 vccd1 _06677_/Y sky130_fd_sc_hd__inv_2
XPHY_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08416_ _08420_/A vssd1 vssd1 vccd1 vccd1 _08416_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09396_ _12454_/Q _10586_/A vssd1 vssd1 vccd1 vccd1 _09396_/X sky130_fd_sc_hd__or2_1
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08347_ _08113_/X _11582_/X _08349_/S vssd1 vssd1 vccd1 vccd1 _12807_/D sky130_fd_sc_hd__mux2_1
XFILLER_149_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_102_wb_clk_i _13235_/CLK vssd1 vssd1 vccd1 vccd1 _13237_/CLK sky130_fd_sc_hd__clkbuf_16
X_08278_ _10411_/A _11610_/S _08278_/C vssd1 vssd1 vccd1 vccd1 _08337_/A sky130_fd_sc_hd__or3_1
XFILLER_192_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07229_ _11568_/X _07218_/X _13103_/Q _07219_/X vssd1 vssd1 vccd1 vccd1 _13103_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10240_ _09595_/Y _10166_/X _10239_/Y _10168_/X vssd1 vssd1 vccd1 vccd1 _10240_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10171_ _10160_/Y _10140_/X _10161_/Y _10141_/X _10170_/X vssd1 vssd1 vccd1 vccd1
+ _10171_/X sky130_fd_sc_hd__o221a_1
XFILLER_160_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput480 _11231_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput491 _11241_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12812_ _12169_/X _12812_/D _08334_/X vssd1 vssd1 vccd1 vccd1 _12812_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_170_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12743_ _12743_/CLK _12743_/D _08591_/X vssd1 vssd1 vccd1 vccd1 _12743_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12679_/CLK _12674_/D _08779_/X vssd1 vssd1 vccd1 vccd1 _12674_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _10495_/X _12992_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11625_/X sky130_fd_sc_hd__mux2_1
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11556_ _12813_/Q _09243_/D _11558_/S vssd1 vssd1 vccd1 vccd1 _11556_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10507_ _12581_/Q _07755_/B _07756_/B vssd1 vssd1 vccd1 vccd1 _10507_/X sky130_fd_sc_hd__a21bo_1
XFILLER_6_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11487_ _10332_/X input356/X _11487_/S vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13226_ _13236_/CLK _13226_/D _06522_/X vssd1 vssd1 vccd1 vccd1 _13226_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10438_ _08187_/X _10439_/C _12816_/Q _10436_/B _10437_/X vssd1 vssd1 vccd1 vccd1
+ _10438_/X sky130_fd_sc_hd__o221a_1
XFILLER_98_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13157_ _13158_/CLK _13157_/D _07055_/X vssd1 vssd1 vccd1 vccd1 _13157_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10369_ _10373_/B vssd1 vssd1 vccd1 vccd1 _10376_/C sky130_fd_sc_hd__inv_2
XFILLER_3_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12108_ _10714_/Y _10715_/Y _12770_/Q vssd1 vssd1 vccd1 vccd1 _12193_/S sky130_fd_sc_hd__mux2_8
X_13088_ _12167_/X _13088_/D _07266_/X vssd1 vssd1 vccd1 vccd1 _13088_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_100_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12039_ _11073_/X _11066_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06600_ _06766_/A vssd1 vssd1 vccd1 vccd1 _06650_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07580_ _12982_/Q _07574_/X _09186_/A _07575_/X _07576_/X vssd1 vssd1 vccd1 vccd1
+ _12982_/D sky130_fd_sc_hd__o221a_1
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06531_ _06531_/A vssd1 vssd1 vccd1 vccd1 _13225_/D sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_0_wb_clk_i clkbuf_opt_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12165_/A0
+ sky130_fd_sc_hd__clkbuf_16
X_09250_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09250_/X sky130_fd_sc_hd__clkbuf_2
X_06462_ _13233_/Q vssd1 vssd1 vccd1 vccd1 _06462_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08201_ _08197_/Y _08113_/X _08198_/Y _10475_/A _08200_/X vssd1 vssd1 vccd1 vccd1
+ _08209_/B sky130_fd_sc_hd__a221o_1
XFILLER_147_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09181_ _09243_/C _09243_/D vssd1 vssd1 vccd1 vccd1 _10529_/A sky130_fd_sc_hd__or2_2
X_06393_ _06382_/X _12214_/X _06375_/X _06392_/X vssd1 vssd1 vccd1 vccd1 _13244_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08132_ _08132_/A _08132_/B _08132_/C _08131_/X vssd1 vssd1 vccd1 vccd1 _08132_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_193_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08063_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08063_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07014_ _07024_/A vssd1 vssd1 vccd1 vccd1 _07014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput208 la_oenb[21] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__buf_1
X_08965_ _08969_/A vssd1 vssd1 vccd1 vccd1 _08965_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_130_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput219 la_oenb[31] vssd1 vssd1 vccd1 vccd1 input219/X sky130_fd_sc_hd__buf_1
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07916_ _07815_/X _11503_/X _07918_/S vssd1 vssd1 vccd1 vccd1 _12914_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08896_ _08883_/X _06311_/Y _08893_/X _12630_/Q vssd1 vssd1 vccd1 vccd1 _12630_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07847_ _12908_/Q vssd1 vssd1 vccd1 vccd1 _10357_/A sky130_fd_sc_hd__inv_2
XFILLER_112_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07778_ _07778_/A _09437_/A vssd1 vssd1 vccd1 vccd1 _07781_/A sky130_fd_sc_hd__or2_2
XFILLER_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09517_ _09502_/X _09505_/Y _09516_/Y vssd1 vssd1 vccd1 vccd1 _09517_/Y sky130_fd_sc_hd__o21ai_1
X_06729_ _06726_/X _06727_/X _12014_/X _06728_/X vssd1 vssd1 vccd1 vccd1 _06729_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _12967_/Q _09440_/X _13003_/Q _09442_/A _09447_/X vssd1 vssd1 vccd1 vccd1
+ _09448_/X sky130_fd_sc_hd__a221o_1
XFILLER_13_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09379_ _12456_/Q vssd1 vssd1 vccd1 vccd1 _09379_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11410_ _12443_/Q _11409_/X _12139_/S vssd1 vssd1 vccd1 vccd1 _11410_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12390_ _12995_/CLK _12390_/D vssd1 vssd1 vccd1 vccd1 _12412_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11341_ vssd1 vssd1 vccd1 vccd1 _11341_/HI _11341_/LO sky130_fd_sc_hd__conb_1
XFILLER_126_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11272_ vssd1 vssd1 vccd1 vccd1 _11272_/HI _11272_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13011_ _12164_/X _13011_/D _07487_/X vssd1 vssd1 vccd1 vccd1 _13011_/Q sky130_fd_sc_hd__dfrtp_4
X_10223_ _10221_/Y _10166_/X _10222_/Y _10168_/X vssd1 vssd1 vccd1 vccd1 _10223_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_70_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12951_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_121_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10154_ _07403_/Y _10090_/X _08475_/Y _10113_/X vssd1 vssd1 vccd1 vccd1 _10154_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10085_ _12774_/Q vssd1 vssd1 vccd1 vccd1 _10085_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10987_ _12540_/Q _12352_/Q _12540_/Q _12352_/Q vssd1 vssd1 vccd1 vccd1 _11000_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_188_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12726_ _12726_/CLK _12726_/D _08636_/X vssd1 vssd1 vccd1 vccd1 _12726_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_71_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ _13264_/CLK _12657_/D _08828_/X vssd1 vssd1 vccd1 vccd1 _12657_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11608_ _10483_/Y _10794_/A _11610_/S vssd1 vssd1 vccd1 vccd1 _11608_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12588_ _12993_/CLK _12588_/D vssd1 vssd1 vccd1 vccd1 _12588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11539_ _12828_/Q _10792_/B _11543_/S vssd1 vssd1 vccd1 vccd1 _11539_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13209_ _13213_/CLK _13209_/D _06687_/X vssd1 vssd1 vccd1 vccd1 _13209_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08750_ _08854_/A vssd1 vssd1 vccd1 vccd1 _08839_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07701_ _12309_/Q vssd1 vssd1 vccd1 vccd1 _07702_/A sky130_fd_sc_hd__inv_2
XFILLER_39_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08681_ _11843_/X _08670_/X _12709_/Q _08671_/X vssd1 vssd1 vccd1 vccd1 _12709_/D
+ sky130_fd_sc_hd__a22o_1
X_07632_ _12947_/Q _12946_/Q _12948_/Q _12953_/Q vssd1 vssd1 vccd1 vccd1 _07650_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_4_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07563_ _07562_/X _07552_/X _12989_/Q _07553_/X _07556_/X vssd1 vssd1 vccd1 vccd1
+ _12989_/D sky130_fd_sc_hd__a221o_1
XFILLER_59_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09302_ _09302_/A _11968_/X vssd1 vssd1 vccd1 vccd1 _09302_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06514_ _06509_/Y _06510_/Y _06511_/Y _06512_/Y vssd1 vssd1 vccd1 vccd1 _06514_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07494_ _07590_/A vssd1 vssd1 vccd1 vccd1 _07775_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09233_ _09233_/A vssd1 vssd1 vccd1 vccd1 _09233_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_142_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06445_ _12767_/Q _12766_/Q vssd1 vssd1 vccd1 vccd1 _06446_/B sky130_fd_sc_hd__and2_1
XFILLER_148_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13219_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_09164_ _09164_/A vssd1 vssd1 vccd1 vccd1 _09164_/X sky130_fd_sc_hd__clkbuf_2
X_06376_ _13249_/Q vssd1 vssd1 vccd1 vccd1 _06376_/X sky130_fd_sc_hd__buf_2
XFILLER_148_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08115_ _12830_/Q vssd1 vssd1 vccd1 vccd1 _10475_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09095_ _12539_/Q _09089_/X _10794_/A _09092_/X vssd1 vssd1 vccd1 vccd1 _12539_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08046_ _12868_/Q _08040_/X _07290_/X _08041_/X vssd1 vssd1 vccd1 vccd1 _12868_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09997_ _08780_/Y _09993_/X _06240_/Y _09972_/X _09991_/X vssd1 vssd1 vccd1 vccd1
+ _09997_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08948_ _12431_/Q _12432_/Q vssd1 vssd1 vccd1 vccd1 _08949_/B sky130_fd_sc_hd__or2_1
XFILLER_130_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08879_ _08877_/X _06271_/Y _12637_/Q _08878_/X vssd1 vssd1 vccd1 vccd1 _12637_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10910_ _10908_/X _10909_/X _10908_/X _10909_/X vssd1 vssd1 vccd1 vccd1 _12340_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11890_ _08925_/A _10628_/Y _12321_/Q vssd1 vssd1 vccd1 vccd1 _11890_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10841_ _12519_/Q vssd1 vssd1 vccd1 vccd1 _10843_/A sky130_fd_sc_hd__inv_2
XFILLER_44_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10772_ _13246_/Q vssd1 vssd1 vccd1 vccd1 _10773_/A sky130_fd_sc_hd__inv_2
XFILLER_73_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _12517_/CLK _12511_/D vssd1 vssd1 vccd1 vccd1 _12511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12442_ _12442_/CLK _12442_/D vssd1 vssd1 vccd1 vccd1 _12442_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12373_ _12376_/CLK _12373_/D vssd1 vssd1 vccd1 vccd1 _12395_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_166_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11324_ vssd1 vssd1 vccd1 vccd1 _11324_/HI _11324_/LO sky130_fd_sc_hd__conb_1
XFILLER_197_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11255_ vssd1 vssd1 vccd1 vccd1 _11255_/HI _11255_/LO sky130_fd_sc_hd__conb_1
XFILLER_153_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10206_ _09914_/Y _10134_/X _10197_/X _10205_/X vssd1 vssd1 vccd1 vccd1 _10206_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_79_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ vssd1 vssd1 vccd1 vccd1 _11186_/HI _11186_/LO sky130_fd_sc_hd__conb_1
XFILLER_80_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10137_ _10137_/A vssd1 vssd1 vccd1 vccd1 _10137_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10068_ _10068_/A _10068_/B _10068_/C _10068_/D vssd1 vssd1 vccd1 vccd1 _10068_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_169_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12709_ _12713_/CLK _12709_/D _08680_/X vssd1 vssd1 vccd1 vccd1 _12709_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06230_ _06245_/A vssd1 vssd1 vccd1 vccd1 _06230_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06161_ _08556_/B _06272_/A vssd1 vssd1 vccd1 vccd1 _06162_/A sky130_fd_sc_hd__or2_1
XFILLER_117_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06092_ _06092_/A vssd1 vssd1 vccd1 vccd1 _06130_/A sky130_fd_sc_hd__inv_2
XFILLER_116_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09920_ _12663_/Q _12611_/Q _06305_/X _09547_/A _09919_/Y vssd1 vssd1 vccd1 vccd1
+ _09920_/X sky130_fd_sc_hd__a221o_1
XFILLER_125_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09851_ _09851_/A _09851_/B vssd1 vssd1 vccd1 vccd1 _09851_/X sky130_fd_sc_hd__or2_1
X_08802_ _08798_/X _08801_/X _06278_/Y _12668_/Q _08567_/X vssd1 vssd1 vccd1 vccd1
+ _12668_/D sky130_fd_sc_hd__a32o_1
XFILLER_86_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09782_ _09782_/A _09782_/B vssd1 vssd1 vccd1 vccd1 _09782_/Y sky130_fd_sc_hd__nor2_1
X_06994_ _07006_/A vssd1 vssd1 vccd1 vccd1 _06994_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08733_ _11822_/X _08592_/A _12688_/Q _08593_/A vssd1 vssd1 vccd1 vccd1 _12688_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08664_ _11850_/X _08654_/X _12716_/Q _08655_/X vssd1 vssd1 vccd1 vccd1 _12716_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07615_ _11615_/X _07610_/X _12970_/Q _07611_/X _07583_/X vssd1 vssd1 vccd1 vccd1
+ _12970_/D sky130_fd_sc_hd__o221a_1
XPHY_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08595_ _08642_/A vssd1 vssd1 vccd1 vccd1 _08606_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ _07778_/A vssd1 vssd1 vccd1 vccd1 _11982_/S sky130_fd_sc_hd__inv_2
XPHY_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07477_ _07477_/A vssd1 vssd1 vccd1 vccd1 _07933_/A sky130_fd_sc_hd__buf_4
XFILLER_195_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09216_ _09216_/A vssd1 vssd1 vccd1 vccd1 _09216_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06428_ _10717_/A vssd1 vssd1 vccd1 vccd1 _10737_/A sky130_fd_sc_hd__buf_2
XFILLER_167_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09147_ _12508_/Q _09147_/B vssd1 vssd1 vccd1 vccd1 _09147_/X sky130_fd_sc_hd__or2_2
XFILLER_148_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06359_ _12234_/X _08504_/A _06356_/X _06358_/X vssd1 vssd1 vccd1 vccd1 _13254_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_163_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09078_ _09247_/A _11703_/S vssd1 vssd1 vccd1 vccd1 _09079_/A sky130_fd_sc_hd__nand2_2
XFILLER_135_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08029_ _12875_/Q _08024_/X _07980_/X _08026_/X vssd1 vssd1 vccd1 vccd1 _12875_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11040_ _10686_/X _10746_/X _06410_/X _07008_/X _10747_/X vssd1 vssd1 vccd1 vccd1
+ _11040_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12991_ _13004_/CLK _12991_/D vssd1 vssd1 vccd1 vccd1 _12991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11942_ _09683_/X _12803_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11942_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11873_ _10246_/X _12814_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11873_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10824_ _12516_/Q vssd1 vssd1 vccd1 vccd1 _10824_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10755_ _10755_/A vssd1 vssd1 vccd1 vccd1 _10755_/X sky130_fd_sc_hd__buf_2
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10686_ _10686_/A vssd1 vssd1 vccd1 vccd1 _10686_/X sky130_fd_sc_hd__buf_2
X_12425_ _12426_/CLK _12425_/D vssd1 vssd1 vccd1 vccd1 _12425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12356_ _12357_/CLK _12356_/D vssd1 vssd1 vccd1 vccd1 _12356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11307_ vssd1 vssd1 vccd1 vccd1 _11307_/HI _11307_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12287_ _12296_/CLK _12287_/D vssd1 vssd1 vccd1 vccd1 _12287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_2_wb_clk_i clkbuf_opt_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _12284_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_45_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11238_ vssd1 vssd1 vccd1 vccd1 _11238_/HI _11238_/LO sky130_fd_sc_hd__conb_1
XFILLER_45_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11169_ vssd1 vssd1 vccd1 vccd1 _11169_/HI _11169_/LO sky130_fd_sc_hd__conb_1
XFILLER_96_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07400_ _07408_/A vssd1 vssd1 vccd1 vccd1 _07400_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08380_ _12795_/Q _08374_/X _07290_/X _08375_/X vssd1 vssd1 vccd1 vccd1 _12795_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07331_ _11446_/X _07321_/X _13070_/Q _07324_/X vssd1 vssd1 vccd1 vccd1 _13070_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07262_ _07266_/A vssd1 vssd1 vccd1 vccd1 _07262_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09001_ _09002_/A _11029_/A vssd1 vssd1 vccd1 vccd1 _12594_/D sky130_fd_sc_hd__or2_1
XFILLER_164_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06213_ _06207_/Y _06022_/X _06163_/X _06212_/X vssd1 vssd1 vccd1 vccd1 _13281_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_117_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07193_ _11515_/X _07160_/A _13114_/Q _07161_/A vssd1 vssd1 vccd1 vccd1 _13114_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06144_ _06144_/A _06144_/B vssd1 vssd1 vccd1 vccd1 _06144_/X sky130_fd_sc_hd__or2_1
XFILLER_133_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06075_ _06075_/A _06075_/B vssd1 vssd1 vccd1 vccd1 _06182_/A sky130_fd_sc_hd__or2_2
XFILLER_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09903_ _12658_/Q vssd1 vssd1 vccd1 vccd1 _09903_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_127_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13286_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09834_ _06508_/Y _09820_/X _06503_/Y _09821_/X vssd1 vssd1 vccd1 vccd1 _09839_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_98_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09765_ _09769_/A _09849_/A _09745_/Y vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__a21oi_2
XFILLER_6_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06977_ _06977_/A _06977_/B vssd1 vssd1 vccd1 vccd1 _06977_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08716_ _08716_/A vssd1 vssd1 vccd1 vccd1 _08716_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09696_ _09696_/A vssd1 vssd1 vccd1 vccd1 _09713_/B sky130_fd_sc_hd__inv_2
XPHY_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08647_ _08653_/A vssd1 vssd1 vccd1 vccd1 _08647_/X sky130_fd_sc_hd__clkbuf_1
XPHY_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08578_ _08593_/A vssd1 vssd1 vccd1 vccd1 _08578_/X sky130_fd_sc_hd__clkbuf_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07529_ _07778_/A _09443_/A vssd1 vssd1 vccd1 vccd1 _07532_/A sky130_fd_sc_hd__or2_2
XPHY_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10540_ _11360_/X _10554_/B vssd1 vssd1 vccd1 vccd1 _10540_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10471_ _08164_/Y _10468_/A _12828_/Q _10472_/C _10437_/X vssd1 vssd1 vccd1 vccd1
+ _10471_/X sky130_fd_sc_hd__o221a_1
XFILLER_194_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12210_ _12209_/X _12625_/Q _12552_/Q vssd1 vssd1 vccd1 vccd1 _12210_/X sky130_fd_sc_hd__mux2_2
X_13190_ _13190_/CLK _13190_/D _06863_/X vssd1 vssd1 vccd1 vccd1 _13190_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_198_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12141_ _12438_/Q _12140_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12141_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12072_ _06535_/A _10704_/Y _12762_/Q vssd1 vssd1 vccd1 vccd1 _12200_/S sky130_fd_sc_hd__mux2_8
XFILLER_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11023_ _12361_/Q vssd1 vssd1 vccd1 vccd1 _11024_/A sky130_fd_sc_hd__inv_2
XFILLER_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12974_ _12974_/CLK _12974_/D vssd1 vssd1 vccd1 vccd1 _12974_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11925_ _10306_/Y _12802_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _11925_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ _10043_/Y _12313_/Q _12312_/Q vssd1 vssd1 vccd1 vccd1 _11856_/X sky130_fd_sc_hd__mux2_2
XFILLER_199_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10807_ _10807_/A vssd1 vssd1 vccd1 vccd1 _10807_/Y sky130_fd_sc_hd__inv_2
XPHY_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11787_ _12130_/X _12481_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11787_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10738_ _10738_/A vssd1 vssd1 vccd1 vccd1 _10738_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10669_ _12431_/Q _09312_/A _12432_/Q vssd1 vssd1 vccd1 vccd1 _10669_/X sky130_fd_sc_hd__o21a_1
XFILLER_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12408_ _12410_/CLK _12408_/D vssd1 vssd1 vccd1 vccd1 _12408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12339_ _12357_/CLK _12339_/D vssd1 vssd1 vccd1 vccd1 _12339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06900_ _12017_/X _06898_/B _06898_/X vssd1 vssd1 vccd1 vccd1 _06900_/X sky130_fd_sc_hd__a21bo_1
X_07880_ _07880_/A _07880_/B _07880_/C _07879_/X vssd1 vssd1 vccd1 vccd1 _07888_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_68_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06831_ _06816_/X _06820_/X _06821_/X vssd1 vssd1 vccd1 vccd1 _06831_/X sky130_fd_sc_hd__a21bo_1
XFILLER_110_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09550_ _09550_/A _09550_/B vssd1 vssd1 vccd1 vccd1 _09550_/Y sky130_fd_sc_hd__nor2_2
X_06762_ _12002_/X _11999_/X _06756_/X _06757_/X _06761_/X vssd1 vssd1 vccd1 vccd1
+ _06762_/X sky130_fd_sc_hd__o32a_2
XFILLER_83_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08501_ _08503_/A vssd1 vssd1 vccd1 vccd1 _08501_/X sky130_fd_sc_hd__clkbuf_1
X_09481_ _13165_/Q vssd1 vssd1 vccd1 vccd1 _09482_/C sky130_fd_sc_hd__inv_2
X_06693_ _12052_/X _06668_/X _12052_/X _06668_/X vssd1 vssd1 vccd1 vccd1 _06694_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ _12775_/Q _08417_/A _07562_/X _08418_/A vssd1 vssd1 vccd1 vccd1 _12775_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08363_ _12802_/Q _08358_/X _07980_/X _08360_/X vssd1 vssd1 vccd1 vccd1 _12802_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07314_ _13074_/Q _07285_/A _07313_/X _07284_/A vssd1 vssd1 vccd1 vccd1 _13074_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08294_ _08353_/S vssd1 vssd1 vccd1 vccd1 _08307_/S sky130_fd_sc_hd__buf_2
XFILLER_192_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07245_ _07251_/A vssd1 vssd1 vccd1 vccd1 _07245_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07176_ _07176_/A vssd1 vssd1 vccd1 vccd1 _07176_/X sky130_fd_sc_hd__buf_2
XFILLER_117_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06127_ _12724_/Q _12692_/Q _06126_/X vssd1 vssd1 vccd1 vccd1 _06176_/A sky130_fd_sc_hd__o21ai_2
XFILLER_105_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06058_ _12736_/Q _12704_/Q _12736_/Q _12704_/Q vssd1 vssd1 vccd1 vccd1 _06060_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09817_ _09817_/A vssd1 vssd1 vccd1 vccd1 _09817_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09748_ _09748_/A _09770_/A _09748_/C vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__or3_4
XFILLER_28_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09679_ _13162_/Q vssd1 vssd1 vccd1 vccd1 _09679_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11709_/X _10634_/Y _11774_/S vssd1 vssd1 vccd1 vccd1 _12419_/D sky130_fd_sc_hd__mux2_1
XPHY_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_95_wb_clk_i _13235_/CLK vssd1 vssd1 vccd1 vccd1 _13183_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12690_ _12695_/CLK _12690_/D _08727_/X vssd1 vssd1 vccd1 vccd1 _12690_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_199_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12442_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _10511_/X _12926_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11641_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _12829_/Q _10792_/A _11578_/S vssd1 vssd1 vccd1 vccd1 _11572_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 io_in[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
X_10523_ _12404_/D _12405_/D vssd1 vssd1 vccd1 vccd1 _10585_/A sky130_fd_sc_hd__or2_1
XPHY_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13242_ _13252_/CLK _13242_/D _06399_/X vssd1 vssd1 vccd1 vccd1 _13242_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10454_ _10454_/A _10454_/B vssd1 vssd1 vccd1 vccd1 _10455_/C sky130_fd_sc_hd__or2_1
XFILLER_6_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13173_ _13177_/CLK _13173_/D _06997_/X vssd1 vssd1 vccd1 vccd1 _13173_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10385_ _12918_/Q _12917_/Q _10385_/C vssd1 vssd1 vccd1 vccd1 _10388_/B sky130_fd_sc_hd__and3_1
X_12124_ _12123_/X _12434_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12124_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12055_ _11053_/X _11047_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12055_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater609 _11819_/S vssd1 vssd1 vccd1 vccd1 _11774_/S sky130_fd_sc_hd__buf_8
X_11006_ _12355_/Q vssd1 vssd1 vccd1 vccd1 _11014_/B sky130_fd_sc_hd__inv_2
XFILLER_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12957_ _12957_/CLK _12957_/D vssd1 vssd1 vccd1 vccd1 _12957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11908_ _12142_/S _12449_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _11908_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12888_/CLK _12888_/D _07989_/X vssd1 vssd1 vccd1 vccd1 _12888_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11839_ _09947_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11839_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07030_ _11034_/A vssd1 vssd1 vccd1 vccd1 _07030_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08981_ _08980_/Y _07637_/Y _07654_/B _12307_/Q _07695_/X vssd1 vssd1 vccd1 vccd1
+ _12602_/D sky130_fd_sc_hd__o311a_1
XFILLER_114_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07932_ _12907_/Q _11496_/X _07932_/S vssd1 vssd1 vccd1 vccd1 _12907_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07863_ _12904_/Q vssd1 vssd1 vccd1 vccd1 _10346_/A sky130_fd_sc_hd__inv_2
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06814_ _12038_/X vssd1 vssd1 vccd1 vccd1 _06815_/B sky130_fd_sc_hd__inv_2
X_09602_ _13188_/Q _09602_/B vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__nand2_1
X_07794_ _13039_/Q vssd1 vssd1 vccd1 vccd1 _07794_/Y sky130_fd_sc_hd__inv_2
X_09533_ _13152_/Q _07737_/A _09532_/Y _09478_/X vssd1 vssd1 vccd1 vccd1 _09533_/X
+ sky130_fd_sc_hd__o22a_1
X_06745_ _06740_/X _06741_/X _06734_/X _06730_/X _06744_/X vssd1 vssd1 vccd1 vccd1
+ _06745_/X sky130_fd_sc_hd__o221a_1
XFILLER_37_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09464_ _12932_/Q _09438_/A _13000_/Q _09451_/X _09463_/X vssd1 vssd1 vccd1 vccd1
+ _09464_/X sky130_fd_sc_hd__a221o_1
XFILLER_58_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06676_ _06690_/A vssd1 vssd1 vccd1 vccd1 _06676_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08415_ _12782_/Q _08401_/X _07993_/X _08403_/X vssd1 vssd1 vccd1 vccd1 _12782_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_196_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09395_ _12406_/D vssd1 vssd1 vccd1 vccd1 _10586_/A sky130_fd_sc_hd__inv_2
XFILLER_145_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08346_ _08352_/A vssd1 vssd1 vccd1 vccd1 _08346_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08277_ _08272_/Y _08274_/X _13078_/Q _08275_/Y _10052_/A vssd1 vssd1 vccd1 vccd1
+ _08278_/C sky130_fd_sc_hd__a221oi_2
XFILLER_192_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07228_ _07236_/A vssd1 vssd1 vccd1 vccd1 _07228_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_180_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_142_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12888_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_106_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07159_ _07167_/A vssd1 vssd1 vccd1 vccd1 _07159_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10170_ _10162_/Y _10163_/X _10164_/Y _10165_/X _10169_/X vssd1 vssd1 vccd1 vccd1
+ _10170_/X sky130_fd_sc_hd__o221a_1
Xoutput470 _11337_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput481 _11232_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_120_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput492 _11242_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_87_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12811_ _12169_/X _12811_/D _08336_/X vssd1 vssd1 vccd1 vccd1 _12811_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_76_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12742_ _12743_/CLK _12742_/D _08596_/X vssd1 vssd1 vccd1 vccd1 _12742_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_103_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12679_/CLK _12673_/D _08783_/X vssd1 vssd1 vccd1 vccd1 _12673_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _10494_/X _12991_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11624_/X sky130_fd_sc_hd__mux2_1
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11555_ _12812_/Q _09183_/A _11558_/S vssd1 vssd1 vccd1 vccd1 _11555_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10506_ _12580_/Q _12579_/Q _07755_/B vssd1 vssd1 vccd1 vccd1 _10506_/X sky130_fd_sc_hd__a21bo_1
XFILLER_171_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11486_ _10330_/Y input355/X _11487_/S vssd1 vssd1 vccd1 vccd1 _11486_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13225_ _13236_/CLK _13225_/D _06525_/X vssd1 vssd1 vccd1 vccd1 _13225_/Q sky130_fd_sc_hd__dfrtp_1
X_10437_ _10459_/A vssd1 vssd1 vccd1 vccd1 _10437_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_152_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13156_ _13156_/CLK _13156_/D _07057_/X vssd1 vssd1 vccd1 vccd1 _13156_/Q sky130_fd_sc_hd__dfrtp_4
X_10368_ _10368_/A _10368_/B _10368_/C _10368_/D vssd1 vssd1 vccd1 vccd1 _10373_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_83_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12107_ _12106_/X _12431_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12107_/X sky130_fd_sc_hd__mux2_1
X_13087_ _12167_/X _13087_/D _07270_/X vssd1 vssd1 vccd1 vccd1 _13087_/Q sky130_fd_sc_hd__dfrtp_4
X_10299_ _12891_/Q vssd1 vssd1 vccd1 vccd1 _10299_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12038_ _11089_/X _11080_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06530_ _06526_/X _06520_/B _06527_/Y _06528_/X _06529_/Y vssd1 vssd1 vccd1 vccd1
+ _06531_/A sky130_fd_sc_hd__o32a_1
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06461_ _06465_/A vssd1 vssd1 vccd1 vccd1 _06461_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08200_ _08198_/Y _12830_/Q _08199_/Y _08117_/X vssd1 vssd1 vccd1 vccd1 _08200_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_178_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09180_ _09180_/A _09180_/B _09180_/C _09180_/D vssd1 vssd1 vccd1 vccd1 _09187_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_18_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06392_ _13244_/Q vssd1 vssd1 vccd1 vccd1 _06392_/X sky130_fd_sc_hd__buf_2
XFILLER_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08131_ _08112_/Y _08113_/X _13137_/Q _10467_/A _08130_/X vssd1 vssd1 vccd1 vccd1
+ _08131_/X sky130_fd_sc_hd__o221a_1
XFILLER_119_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08062_ _12861_/Q _08040_/A _07313_/X _08041_/A vssd1 vssd1 vccd1 vccd1 _12861_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07013_ _06528_/X _07003_/Y _07012_/X _06435_/X _13171_/Q vssd1 vssd1 vccd1 vccd1
+ _13171_/D sky130_fd_sc_hd__a32o_1
XFILLER_162_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput209 la_oenb[22] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__buf_1
X_08964_ _08969_/A vssd1 vssd1 vccd1 vccd1 _08964_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07915_ _07917_/A vssd1 vssd1 vccd1 vccd1 _07915_/X sky130_fd_sc_hd__clkbuf_1
X_08895_ _08897_/A vssd1 vssd1 vccd1 vccd1 _08895_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07846_ _12898_/Q vssd1 vssd1 vccd1 vccd1 _10331_/A sky130_fd_sc_hd__inv_2
XFILLER_57_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07777_ _09441_/A _10527_/B _09982_/B vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__or3_4
XFILLER_140_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06728_ _06726_/X _06727_/X _06726_/X _06727_/X vssd1 vssd1 vccd1 vccd1 _06728_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09516_ _09521_/B vssd1 vssd1 vccd1 vccd1 _09516_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _12603_/Q _07519_/B _12995_/Q _09451_/A vssd1 vssd1 vccd1 vccd1 _09447_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06659_ _13213_/Q vssd1 vssd1 vccd1 vccd1 _06659_/Y sky130_fd_sc_hd__inv_2
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ _09366_/Y _12399_/Q _09374_/Y _12411_/Q _09377_/X vssd1 vssd1 vccd1 vccd1
+ _09382_/C sky130_fd_sc_hd__o221a_1
XFILLER_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08329_ _12815_/Q _11590_/X _08335_/S vssd1 vssd1 vccd1 vccd1 _12815_/D sky130_fd_sc_hd__mux2_1
XFILLER_165_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11340_ vssd1 vssd1 vccd1 vccd1 _11340_/HI _11340_/LO sky130_fd_sc_hd__conb_1
XFILLER_181_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11271_ vssd1 vssd1 vccd1 vccd1 _11271_/HI _11271_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13010_ _12164_/X _13010_/D _07489_/X vssd1 vssd1 vccd1 vccd1 _13010_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10222_ _12647_/Q vssd1 vssd1 vccd1 vccd1 _10222_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _08239_/Y _10151_/X _10152_/X vssd1 vssd1 vccd1 vccd1 _10153_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_160_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10084_ _12753_/Q vssd1 vssd1 vccd1 vccd1 _10084_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10986_ _10983_/Y _10985_/A _11000_/B _10985_/Y vssd1 vssd1 vccd1 vccd1 _12351_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12725_ _12725_/CLK _12725_/D _08638_/X vssd1 vssd1 vccd1 vccd1 _12725_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_128_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ _13264_/CLK _12656_/D _08830_/X vssd1 vssd1 vccd1 vccd1 _12656_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11607_ _10481_/X _10794_/B _11610_/S vssd1 vssd1 vccd1 vccd1 _11607_/X sky130_fd_sc_hd__mux2_1
X_12587_ _12993_/CLK _12587_/D vssd1 vssd1 vccd1 vccd1 _12587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11538_ _12827_/Q _09179_/C _11543_/S vssd1 vssd1 vccd1 vccd1 _11538_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11469_ _12912_/Q _09180_/C _11469_/S vssd1 vssd1 vccd1 vccd1 _11469_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13208_ _13208_/CLK _13208_/D _06690_/X vssd1 vssd1 vccd1 vccd1 _13208_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13139_ _12168_/X _13139_/D _07129_/X vssd1 vssd1 vccd1 vccd1 _13139_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07700_ _12960_/Q _07694_/X _12959_/Q _07698_/X _07695_/X vssd1 vssd1 vccd1 vccd1
+ _12960_/D sky130_fd_sc_hd__o221a_1
X_08680_ _08684_/A vssd1 vssd1 vccd1 vccd1 _08680_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07631_ _07678_/C vssd1 vssd1 vccd1 vccd1 _07631_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07562_ _07562_/A vssd1 vssd1 vccd1 vccd1 _07562_/X sky130_fd_sc_hd__buf_4
XFILLER_179_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09301_ _12942_/Q _12941_/Q _09986_/B vssd1 vssd1 vccd1 vccd1 _09301_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_80_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06513_ _12162_/X _12161_/X _06511_/Y _06512_/Y vssd1 vssd1 vccd1 vccd1 _06549_/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_146_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07493_ _11450_/X _07459_/A _13009_/Q _07460_/A vssd1 vssd1 vccd1 vccd1 _13009_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09232_ _09232_/A vssd1 vssd1 vccd1 vccd1 _09233_/A sky130_fd_sc_hd__inv_2
XFILLER_142_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06444_ _06444_/A _06444_/B vssd1 vssd1 vccd1 vccd1 _06444_/Y sky130_fd_sc_hd__nor2_2
XFILLER_142_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09163_ _09163_/A vssd1 vssd1 vccd1 vccd1 _09163_/X sky130_fd_sc_hd__clkbuf_2
X_06375_ _06396_/A vssd1 vssd1 vccd1 vccd1 _06375_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08114_ _13140_/Q vssd1 vssd1 vccd1 vccd1 _08114_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09094_ _12540_/Q _09089_/X _10793_/B _09092_/X vssd1 vssd1 vccd1 vccd1 _12540_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08045_ _08051_/A vssd1 vssd1 vccd1 vccd1 _08045_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09996_ _08784_/Y _09993_/X _06246_/Y _09972_/X _09991_/X vssd1 vssd1 vccd1 vccd1
+ _09996_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_130_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08947_ _12429_/Q _12430_/Q vssd1 vssd1 vccd1 vccd1 _09312_/A sky130_fd_sc_hd__or2_2
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08878_ _12612_/Q vssd1 vssd1 vccd1 vccd1 _08878_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07829_ _12907_/Q vssd1 vssd1 vccd1 vccd1 _10357_/B sky130_fd_sc_hd__inv_2
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10840_ _10836_/Y _10864_/A _10836_/Y _10864_/A vssd1 vssd1 vccd1 vccd1 _12330_/D
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10771_ _10767_/X _10768_/X _06383_/X _10769_/X _10770_/X vssd1 vssd1 vccd1 vccd1
+ _10771_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12510_ _12517_/CLK _12510_/D vssd1 vssd1 vccd1 vccd1 _12510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ _12441_/CLK _12441_/D vssd1 vssd1 vccd1 vccd1 _12441_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12372_ _12376_/CLK _12372_/D vssd1 vssd1 vccd1 vccd1 _12372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11323_ vssd1 vssd1 vccd1 vccd1 _11323_/HI _11323_/LO sky130_fd_sc_hd__conb_1
XFILLER_154_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11254_ vssd1 vssd1 vccd1 vccd1 _11254_/HI _11254_/LO sky130_fd_sc_hd__conb_1
XFILLER_107_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10205_ _10198_/Y _10140_/X _10199_/Y _10141_/X _10204_/X vssd1 vssd1 vccd1 vccd1
+ _10205_/X sky130_fd_sc_hd__o221a_1
XFILLER_192_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11185_ vssd1 vssd1 vccd1 vccd1 _11185_/HI _11185_/LO sky130_fd_sc_hd__conb_1
X_10136_ _12850_/Q vssd1 vssd1 vccd1 vccd1 _10136_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10067_ _10063_/Y _09999_/A _10064_/Y _10033_/X _10066_/X vssd1 vssd1 vccd1 vccd1
+ _10068_/D sky130_fd_sc_hd__o221a_1
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10969_ _12537_/Q vssd1 vssd1 vccd1 vccd1 _10969_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12708_ _12713_/CLK _12708_/D _08682_/X vssd1 vssd1 vccd1 vccd1 _12708_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12639_ _12870_/CLK _12639_/D _08871_/X vssd1 vssd1 vccd1 vccd1 _12639_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06160_ _12608_/Q vssd1 vssd1 vccd1 vccd1 _08556_/B sky130_fd_sc_hd__inv_2
XFILLER_106_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06091_ _06091_/A _06091_/B vssd1 vssd1 vccd1 vccd1 _06092_/A sky130_fd_sc_hd__or2_1
XFILLER_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09850_ _09827_/Y _09868_/A _09839_/X vssd1 vssd1 vccd1 vccd1 _09881_/A sky130_fd_sc_hd__o21a_1
XFILLER_98_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08801_ _08817_/A vssd1 vssd1 vccd1 vccd1 _08801_/X sky130_fd_sc_hd__clkbuf_2
X_09781_ _09779_/A _09779_/B _09780_/Y vssd1 vssd1 vccd1 vccd1 _09782_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06993_ _06457_/X _09552_/B _06459_/X _06992_/X vssd1 vssd1 vccd1 vccd1 _13175_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_86_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08732_ _08747_/A vssd1 vssd1 vccd1 vccd1 _08732_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08663_ _08669_/A vssd1 vssd1 vccd1 vccd1 _08663_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07614_ _11616_/X _07610_/X _12971_/Q _07611_/X _07583_/X vssd1 vssd1 vccd1 vccd1
+ _12971_/D sky130_fd_sc_hd__o221a_1
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _11952_/X _08592_/X _12743_/Q _08593_/X vssd1 vssd1 vccd1 vccd1 _12743_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07545_ _09185_/A vssd1 vssd1 vccd1 vccd1 _07545_/X sky130_fd_sc_hd__buf_4
XPHY_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07476_ _11457_/X _07474_/X _13016_/Q _07475_/X vssd1 vssd1 vccd1 vccd1 _13016_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09215_ _09215_/A vssd1 vssd1 vccd1 vccd1 _09215_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06427_ _06427_/A vssd1 vssd1 vccd1 vccd1 _06427_/X sky130_fd_sc_hd__buf_2
XFILLER_195_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09146_ _12507_/Q _09146_/B vssd1 vssd1 vccd1 vccd1 _09147_/B sky130_fd_sc_hd__or2_1
XFILLER_154_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06358_ _06396_/A vssd1 vssd1 vccd1 vccd1 _06358_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09077_ _09076_/Y _09180_/B _09180_/A vssd1 vssd1 vccd1 vccd1 _11703_/S sky130_fd_sc_hd__nand3b_4
XFILLER_163_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06289_ _06082_/Y _06083_/Y _06132_/C _06180_/B vssd1 vssd1 vccd1 vccd1 _06289_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_151_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_49_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12547_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08028_ _08036_/A vssd1 vssd1 vccd1 vccd1 _08028_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_200_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09979_ _09975_/Y _10137_/A _09977_/Y _10140_/A vssd1 vssd1 vccd1 vccd1 _09979_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12990_ _12992_/CLK _12990_/D vssd1 vssd1 vccd1 vccd1 _12990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11941_ _09662_/Y _12802_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11941_/X sky130_fd_sc_hd__mux2_2
XFILLER_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11872_ _10230_/X _12813_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11872_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10823_ _12515_/Q _12327_/Q _10822_/X vssd1 vssd1 vccd1 vccd1 _10828_/B sky130_fd_sc_hd__o21a_1
XFILLER_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ _13250_/Q vssd1 vssd1 vccd1 vccd1 _10755_/A sky130_fd_sc_hd__inv_2
XFILLER_185_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10685_ _13239_/Q vssd1 vssd1 vccd1 vccd1 _10686_/A sky130_fd_sc_hd__inv_2
XFILLER_185_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12424_ _12620_/CLK _12424_/D vssd1 vssd1 vccd1 vccd1 _12424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12355_ _12751_/CLK _12355_/D vssd1 vssd1 vccd1 vccd1 _12355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ vssd1 vssd1 vccd1 vccd1 _11306_/HI _11306_/LO sky130_fd_sc_hd__conb_1
XFILLER_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12286_ _12296_/CLK _12286_/D vssd1 vssd1 vccd1 vccd1 _12286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11237_ vssd1 vssd1 vccd1 vccd1 _11237_/HI _11237_/LO sky130_fd_sc_hd__conb_1
XFILLER_49_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11168_ vssd1 vssd1 vccd1 vccd1 _11168_/HI _11168_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10119_ _12642_/Q vssd1 vssd1 vccd1 vccd1 _10119_/Y sky130_fd_sc_hd__inv_2
X_11099_ _11099_/A vssd1 vssd1 vccd1 vccd1 _11099_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07330_ _07330_/A vssd1 vssd1 vccd1 vccd1 _07330_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07261_ _11555_/X _07248_/X _13090_/Q _07249_/X vssd1 vssd1 vccd1 vccd1 _13090_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09000_ _12936_/Q _12934_/Q _12935_/Q _08999_/X _07522_/A vssd1 vssd1 vccd1 vccd1
+ _12595_/D sky130_fd_sc_hd__a221o_1
X_06212_ _06037_/A _06211_/Y _06037_/A _06211_/Y vssd1 vssd1 vccd1 vccd1 _06212_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_164_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07192_ _07206_/A vssd1 vssd1 vccd1 vccd1 _07192_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06143_ _06172_/B _06140_/X _06142_/Y vssd1 vssd1 vccd1 vccd1 _06144_/B sky130_fd_sc_hd__o21a_1
XFILLER_118_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06074_ _12731_/Q _12699_/Q _06072_/Y _06073_/Y vssd1 vssd1 vccd1 vccd1 _06075_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09902_ _09900_/Y _09897_/X _06336_/A _09892_/X _09901_/X vssd1 vssd1 vccd1 vccd1
+ _09902_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09833_ _09701_/X _09831_/Y _09842_/A _09682_/X vssd1 vssd1 vccd1 vccd1 _09833_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_101_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09764_ _09769_/B vssd1 vssd1 vccd1 vccd1 _09764_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06976_ _07006_/A vssd1 vssd1 vccd1 vccd1 _06976_/X sky130_fd_sc_hd__clkbuf_1
X_08715_ _08715_/A vssd1 vssd1 vccd1 vccd1 _08715_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09695_ _09669_/A _09694_/A _09669_/Y _09694_/Y vssd1 vssd1 vccd1 vccd1 _09696_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _11932_/X _08639_/X _12723_/Q _08640_/X vssd1 vssd1 vccd1 vccd1 _12723_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08577_ _08716_/A vssd1 vssd1 vccd1 vccd1 _08593_/A sky130_fd_sc_hd__buf_2
XFILLER_81_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07528_ _10527_/A _09435_/B _09982_/B vssd1 vssd1 vccd1 vccd1 _09443_/A sky130_fd_sc_hd__or3_4
XPHY_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07459_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07459_/X sky130_fd_sc_hd__buf_2
XPHY_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10470_ _10474_/A _10472_/C _10470_/C vssd1 vssd1 vccd1 vccd1 _10470_/Y sky130_fd_sc_hd__nor3_1
XFILLER_182_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09129_ _12513_/Q _09123_/X _07562_/X _09124_/X vssd1 vssd1 vccd1 vccd1 _12513_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12140_ _12139_/X _12438_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12140_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12071_ _12070_/X _12445_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12071_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ _12360_/Q _11021_/B _11024_/B vssd1 vssd1 vccd1 vccd1 _12360_/D sky130_fd_sc_hd__o21a_1
XFILLER_150_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12973_ _12973_/CLK _12973_/D vssd1 vssd1 vccd1 vccd1 _12973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11924_ _10291_/Y _12801_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _11924_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _10053_/X _12804_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11855_/X sky130_fd_sc_hd__mux2_1
XPHY_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ _10806_/A vssd1 vssd1 vccd1 vccd1 _10806_/Y sky130_fd_sc_hd__inv_2
XPHY_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11786_ _11785_/X _12120_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12436_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10737_ _10737_/A vssd1 vssd1 vccd1 vccd1 _10737_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ _12431_/Q _09312_/A _12431_/Q _09312_/A vssd1 vssd1 vccd1 vccd1 _10668_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12407_ _12455_/CLK _12407_/D vssd1 vssd1 vccd1 vccd1 _12407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _10599_/A _10599_/B vssd1 vssd1 vccd1 vccd1 _10603_/B sky130_fd_sc_hd__or2_2
XFILLER_114_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12338_ _12344_/CLK _12338_/D vssd1 vssd1 vccd1 vccd1 _12338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12269_ _10094_/Y _12895_/Q _11859_/X _11860_/X _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12285_/D sky130_fd_sc_hd__mux4_2
XFILLER_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06830_ _13195_/Q vssd1 vssd1 vccd1 vccd1 _06830_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06761_ _06758_/X _06759_/X _12004_/X _06760_/X vssd1 vssd1 vccd1 vccd1 _06761_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08500_ _06403_/X _12264_/X _08499_/X _12769_/Q vssd1 vssd1 vccd1 vccd1 _12769_/D
+ sky130_fd_sc_hd__o22a_1
X_06692_ _11988_/X _11985_/X _11991_/X _06691_/X vssd1 vssd1 vccd1 vccd1 _06694_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09480_ _09471_/X _09474_/X _09479_/X vssd1 vssd1 vccd1 vccd1 _09480_/X sky130_fd_sc_hd__a21bo_1
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08431_ _08433_/A vssd1 vssd1 vccd1 vccd1 _08431_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08362_ _08370_/A vssd1 vssd1 vccd1 vccd1 _08362_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07313_ _07568_/A vssd1 vssd1 vccd1 vccd1 _07313_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08293_ _08296_/A vssd1 vssd1 vccd1 vccd1 _08293_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07244_ _11562_/X _07233_/X _13097_/Q _07234_/X vssd1 vssd1 vccd1 vccd1 _13097_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07175_ _07183_/A vssd1 vssd1 vccd1 vccd1 _07175_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06126_ _12724_/Q _12692_/Q _12723_/Q _12691_/Q vssd1 vssd1 vccd1 vccd1 _06126_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06057_ _06209_/A _06172_/A vssd1 vssd1 vccd1 vccd1 _06144_/A sky130_fd_sc_hd__or2_1
XFILLER_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09816_ _09800_/A _09800_/B _09808_/X vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__o21ai_1
XFILLER_143_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09747_ _09747_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09770_/A sky130_fd_sc_hd__nand2_1
XFILLER_74_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06959_ _11886_/X vssd1 vssd1 vccd1 vccd1 _06960_/B sky130_fd_sc_hd__inv_2
XFILLER_28_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09678_ _09713_/A _09748_/C vssd1 vssd1 vccd1 vccd1 _09678_/Y sky130_fd_sc_hd__nand2_1
XPHY_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08629_ _11939_/X _08624_/X _12730_/Q _08625_/X vssd1 vssd1 vccd1 vccd1 _12730_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _10510_/X _12993_/Q _11648_/S vssd1 vssd1 vccd1 vccd1 _11640_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ _12828_/Q _10792_/B _11578_/S vssd1 vssd1 vccd1 vccd1 _11571_/X sky130_fd_sc_hd__mux2_1
XPHY_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_64_wb_clk_i _12960_/CLK vssd1 vssd1 vccd1 vccd1 _12939_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10522_ _10526_/A vssd1 vssd1 vccd1 vccd1 _10522_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13241_ _13241_/CLK _13241_/D _06402_/X vssd1 vssd1 vccd1 vccd1 _13241_/Q sky130_fd_sc_hd__dfrtp_2
X_10453_ _10454_/B _10450_/A _12822_/Q _10452_/B _10437_/X vssd1 vssd1 vccd1 vccd1
+ _10453_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10384_ _07868_/Y _10381_/A _12917_/Q _10385_/C _10350_/X vssd1 vssd1 vccd1 vccd1
+ _10384_/X sky130_fd_sc_hd__o221a_1
X_13172_ _13177_/CLK _13172_/D _07006_/X vssd1 vssd1 vccd1 vccd1 _13172_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_184_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12123_ _12434_/Q _12122_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12123_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12054_ _11056_/X _11048_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _12054_/X sky130_fd_sc_hd__mux2_2
XFILLER_104_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11005_ _11014_/A _11014_/D _11004_/Y vssd1 vssd1 vccd1 vccd1 _12354_/D sky130_fd_sc_hd__a21oi_1
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12956_ _12957_/CLK _12956_/D vssd1 vssd1 vccd1 vccd1 _12956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11907_ _10650_/Y _10651_/X _12321_/Q vssd1 vssd1 vccd1 vccd1 _11907_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _12888_/CLK _12887_/D _07992_/X vssd1 vssd1 vccd1 vccd1 _12887_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11838_ _09946_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11838_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11769_ _12111_/X _11768_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11769_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08980_ _08980_/A vssd1 vssd1 vccd1 vccd1 _08980_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07931_ _07931_/A vssd1 vssd1 vccd1 vccd1 _07931_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07862_ _12911_/Q vssd1 vssd1 vccd1 vccd1 _10367_/B sky130_fd_sc_hd__inv_2
XFILLER_3_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09601_ _06891_/Y _09600_/Y _13187_/Q _09600_/A vssd1 vssd1 vccd1 vccd1 _09602_/B
+ sky130_fd_sc_hd__o22a_1
X_06813_ _06813_/A _06813_/B vssd1 vssd1 vccd1 vccd1 _06813_/X sky130_fd_sc_hd__or2_1
XFILLER_83_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07793_ _07903_/A vssd1 vssd1 vccd1 vccd1 _07793_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09532_ _12866_/Q vssd1 vssd1 vccd1 vccd1 _09532_/Y sky130_fd_sc_hd__inv_2
X_06744_ _06748_/A _06748_/B vssd1 vssd1 vccd1 vccd1 _06744_/X sky130_fd_sc_hd__or2_1
XFILLER_3_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09463_ _12972_/Q _09440_/A _12599_/Q _07519_/B vssd1 vssd1 vccd1 vccd1 _09463_/X
+ sky130_fd_sc_hd__a22o_1
X_06675_ _06663_/X _06671_/Y _06680_/A _06436_/X _13212_/Q vssd1 vssd1 vccd1 vccd1
+ _13212_/D sky130_fd_sc_hd__o32a_1
XFILLER_52_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08414_ _08420_/A vssd1 vssd1 vccd1 vccd1 _08414_/X sky130_fd_sc_hd__clkbuf_1
X_09394_ _09394_/A vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_196_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08345_ _12808_/Q _11583_/X _08349_/S vssd1 vssd1 vccd1 vccd1 _12808_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08276_ _13074_/Q vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__inv_2
XFILLER_20_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07227_ _11569_/X _07218_/X _13104_/Q _07219_/X vssd1 vssd1 vccd1 vccd1 _13104_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07158_ _11529_/X _07145_/X _13128_/Q _07146_/X vssd1 vssd1 vccd1 vccd1 _13128_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06109_ _12722_/Q _12690_/Q _12721_/Q _12689_/Q vssd1 vssd1 vccd1 vccd1 _06109_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07089_ _11969_/S vssd1 vssd1 vccd1 vccd1 _09984_/A sky130_fd_sc_hd__inv_2
XFILLER_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput460 _11328_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput471 _11338_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__clkbuf_2
Xoutput482 _11233_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput493 _11243_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__clkbuf_2
XFILLER_59_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_111_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 _12749_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12810_ _12169_/X _12810_/D _08339_/X vssd1 vssd1 vccd1 vccd1 _12810_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12741_ _12743_/CLK _12741_/D _08598_/X vssd1 vssd1 vccd1 vccd1 _12741_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12682_/CLK _12672_/D _08786_/X vssd1 vssd1 vccd1 vccd1 _12672_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_42_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _10493_/X _12990_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11623_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11554_ _12811_/Q _09185_/A _11558_/S vssd1 vssd1 vccd1 vccd1 _11554_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10505_ _12579_/Q vssd1 vssd1 vccd1 vccd1 _10505_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11485_ _10327_/X _09186_/B _11487_/S vssd1 vssd1 vccd1 vccd1 _11485_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13224_ _13236_/CLK _13224_/D _06532_/X vssd1 vssd1 vccd1 vccd1 _13224_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10436_ _10458_/A _10436_/B _10436_/C vssd1 vssd1 vccd1 vccd1 _10436_/Y sky130_fd_sc_hd__nor3_2
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13155_ _13156_/CLK _13155_/D _07061_/X vssd1 vssd1 vccd1 vccd1 _13155_/Q sky130_fd_sc_hd__dfrtp_1
X_10367_ _10367_/A _10367_/B vssd1 vssd1 vccd1 vccd1 _10368_/C sky130_fd_sc_hd__or2_1
XFILLER_98_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12106_ _12105_/X _12431_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12106_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10298_ _12786_/Q vssd1 vssd1 vccd1 vccd1 _10298_/Y sky130_fd_sc_hd__inv_2
X_13086_ _12167_/X _13086_/D _07272_/X vssd1 vssd1 vccd1 vccd1 _13086_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12037_ _11095_/X _11090_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12037_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12939_ _12939_/CLK _12939_/D vssd1 vssd1 vccd1 vccd1 _12939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06460_ _06457_/X _06453_/Y _06458_/X _06459_/X _13234_/Q vssd1 vssd1 vccd1 vccd1
+ _13234_/D sky130_fd_sc_hd__a32o_1
XFILLER_22_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06391_ _06391_/A vssd1 vssd1 vccd1 vccd1 _06391_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08130_ _08127_/Y _08128_/X _08129_/Y _12813_/Q vssd1 vssd1 vccd1 vccd1 _08130_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_193_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08061_ _08070_/A vssd1 vssd1 vccd1 vccd1 _08061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_147_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07012_ _07012_/A _07012_/B vssd1 vssd1 vccd1 vccd1 _07012_/X sky130_fd_sc_hd__or2_1
XFILLER_128_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08963_ _08963_/A vssd1 vssd1 vccd1 vccd1 _08969_/A sky130_fd_sc_hd__clkbuf_4
X_07914_ _12915_/Q _11504_/X _07918_/S vssd1 vssd1 vccd1 vccd1 _12915_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08894_ _08883_/X _06305_/A _08893_/X _12631_/Q vssd1 vssd1 vccd1 vccd1 _12631_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07845_ _12903_/Q vssd1 vssd1 vccd1 vccd1 _10346_/B sky130_fd_sc_hd__inv_2
XFILLER_110_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07776_ _12576_/Q _07768_/A _12934_/Q _07769_/X _07775_/X vssd1 vssd1 vccd1 vccd1
+ _12934_/D sky130_fd_sc_hd__a221o_1
XFILLER_72_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09515_ _09500_/A _09500_/B _09514_/A _09500_/Y _09514_/Y vssd1 vssd1 vccd1 vccd1
+ _09521_/B sky130_fd_sc_hd__o32a_1
XFILLER_83_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06727_ _12009_/X _12035_/X _12009_/X _12035_/X vssd1 vssd1 vccd1 vccd1 _06727_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _12978_/Q _09436_/X _12926_/Q _09438_/X _09445_/X vssd1 vssd1 vccd1 vccd1
+ _09446_/X sky130_fd_sc_hd__a221o_1
XFILLER_80_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ _06658_/A vssd1 vssd1 vccd1 vccd1 _06658_/X sky130_fd_sc_hd__buf_2
XFILLER_40_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09377_ _09375_/Y _12407_/Q _12455_/Q _09376_/Y vssd1 vssd1 vccd1 vccd1 _09377_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_12_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06589_ _12200_/X _06587_/B _06587_/X vssd1 vssd1 vccd1 vccd1 _06589_/X sky130_fd_sc_hd__a21bo_1
XFILLER_178_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08328_ _08339_/A vssd1 vssd1 vccd1 vccd1 _08328_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_138_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08259_ _08284_/A vssd1 vssd1 vccd1 vccd1 _08282_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11270_ vssd1 vssd1 vccd1 vccd1 _11270_/HI _11270_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ _13156_/Q vssd1 vssd1 vccd1 vccd1 _10221_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10152_ _07084_/Y _10090_/X _08165_/Y _10113_/X vssd1 vssd1 vccd1 vccd1 _10152_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10083_ _13257_/Q vssd1 vssd1 vccd1 vccd1 _10083_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10985_ _10985_/A vssd1 vssd1 vccd1 vccd1 _10985_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12724_ _13162_/CLK _12724_/D _08643_/X vssd1 vssd1 vccd1 vccd1 _12724_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ _13268_/CLK _12655_/D _08832_/X vssd1 vssd1 vccd1 vccd1 _12655_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ _10479_/Y _10794_/C _11610_/S vssd1 vssd1 vccd1 vccd1 _11606_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12586_ _12586_/CLK _12586_/D vssd1 vssd1 vccd1 vccd1 _12586_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11537_ _12826_/Q _09179_/D _11543_/S vssd1 vssd1 vccd1 vccd1 _11537_/X sky130_fd_sc_hd__mux2_1
XPHY_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11468_ _12911_/Q _09180_/D _11469_/S vssd1 vssd1 vccd1 vccd1 _11468_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13207_ _13208_/CLK _13207_/D _06709_/X vssd1 vssd1 vccd1 vccd1 _13207_/Q sky130_fd_sc_hd__dfrtp_1
X_10419_ _12809_/Q _10416_/Y _10420_/B _10407_/X vssd1 vssd1 vccd1 vccd1 _10419_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11399_ _10621_/Y _12413_/D _11889_/S vssd1 vssd1 vccd1 vccd1 _11399_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13138_ _12168_/X _13138_/D _07133_/X vssd1 vssd1 vccd1 vccd1 _13138_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_97_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13069_ _12165_/X _13069_/D _07333_/X vssd1 vssd1 vccd1 vccd1 _13069_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07630_ _12948_/Q _07670_/C vssd1 vssd1 vccd1 vccd1 _07678_/C sky130_fd_sc_hd__or2_2
XFILLER_38_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07561_ _07560_/X _07552_/X _12990_/Q _07553_/X _07556_/X vssd1 vssd1 vccd1 vccd1
+ _12990_/D sky130_fd_sc_hd__a221o_1
XFILLER_59_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09300_ _09982_/D _11969_/X vssd1 vssd1 vccd1 vccd1 _09300_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06512_ _12161_/X vssd1 vssd1 vccd1 vccd1 _06512_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07492_ _07749_/A vssd1 vssd1 vccd1 vccd1 _07492_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09231_ _09232_/A vssd1 vssd1 vccd1 vccd1 _09231_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06443_ _12194_/X vssd1 vssd1 vccd1 vccd1 _06444_/B sky130_fd_sc_hd__inv_2
XFILLER_107_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09162_ _11629_/X _09154_/X _12504_/Q _09156_/X vssd1 vssd1 vccd1 vccd1 _12504_/D
+ sky130_fd_sc_hd__a22o_1
X_06374_ _06391_/A vssd1 vssd1 vccd1 vccd1 _06374_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08113_ _12807_/Q vssd1 vssd1 vccd1 vccd1 _08113_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09093_ _12541_/Q _09089_/X _10793_/A _09092_/X vssd1 vssd1 vccd1 vccd1 _12541_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08044_ _12869_/Q _08040_/X _07287_/X _08041_/X vssd1 vssd1 vccd1 vccd1 _12869_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09995_ _08787_/Y _09993_/X _06252_/Y _09972_/X _09991_/X vssd1 vssd1 vccd1 vccd1
+ _09995_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_153_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08946_ _12447_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _08953_/B sky130_fd_sc_hd__or2_1
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08877_ _08898_/A vssd1 vssd1 vccd1 vccd1 _08877_/X sky130_fd_sc_hd__buf_2
XFILLER_151_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07828_ _12910_/Q vssd1 vssd1 vccd1 vccd1 _10368_/A sky130_fd_sc_hd__inv_2
XFILLER_151_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07759_ _12585_/Q _07759_/B vssd1 vssd1 vccd1 vccd1 _07760_/B sky130_fd_sc_hd__or2_1
XFILLER_53_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10770_ _12132_/X vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09429_ _12544_/Q _10619_/A _12543_/Q _10611_/B vssd1 vssd1 vccd1 vccd1 _09429_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12440_ _12485_/CLK _12440_/D vssd1 vssd1 vccd1 vccd1 _12440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12371_ _12426_/CLK _12371_/D vssd1 vssd1 vccd1 vccd1 _12371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11322_ vssd1 vssd1 vccd1 vccd1 _11322_/HI _11322_/LO sky130_fd_sc_hd__conb_1
XFILLER_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11253_ vssd1 vssd1 vccd1 vccd1 _11253_/HI _11253_/LO sky130_fd_sc_hd__conb_1
XFILLER_109_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10204_ _10200_/Y _10163_/X _10201_/Y _10165_/X _10203_/X vssd1 vssd1 vccd1 vccd1
+ _10204_/X sky130_fd_sc_hd__o221a_1
XFILLER_79_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11184_ vssd1 vssd1 vccd1 vccd1 _11184_/HI _11184_/LO sky130_fd_sc_hd__conb_1
XFILLER_192_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10135_ _13260_/Q vssd1 vssd1 vccd1 vccd1 _10135_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10066_ _10792_/D _10151_/A _08546_/Y _10065_/Y _10038_/X vssd1 vssd1 vccd1 vccd1
+ _10066_/X sky130_fd_sc_hd__o32a_1
XFILLER_76_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10968_ _10976_/A _10967_/X _10976_/A _10967_/X vssd1 vssd1 vccd1 vccd1 _12348_/D
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_31_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _12707_/CLK _12707_/D _08684_/X vssd1 vssd1 vccd1 vccd1 _12707_/Q sky130_fd_sc_hd__dfrtp_4
X_10899_ _12339_/Q vssd1 vssd1 vccd1 vccd1 _10900_/B sky130_fd_sc_hd__inv_2
XFILLER_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12638_ _12870_/CLK _12638_/D _08873_/X vssd1 vssd1 vccd1 vccd1 _12638_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12569_ _12570_/CLK _12569_/D vssd1 vssd1 vccd1 vccd1 _12569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06090_ _06090_/A vssd1 vssd1 vccd1 vccd1 _06091_/B sky130_fd_sc_hd__inv_2
XFILLER_89_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08800_ _08807_/A vssd1 vssd1 vccd1 vccd1 _08800_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_140_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09780_ _09780_/A vssd1 vssd1 vccd1 vccd1 _09780_/Y sky130_fd_sc_hd__inv_2
X_06992_ _06987_/Y _11882_/X _06991_/Y vssd1 vssd1 vccd1 vccd1 _06992_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08731_ _08731_/A vssd1 vssd1 vccd1 vccd1 _08747_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08662_ _11851_/X _08654_/X _12717_/Q _08655_/X vssd1 vssd1 vccd1 vccd1 _12717_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07613_ _11617_/X _07610_/X _12972_/Q _07611_/X _07583_/X vssd1 vssd1 vccd1 vccd1
+ _12972_/D sky130_fd_sc_hd__o221a_1
XFILLER_199_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08593_ _08593_/A vssd1 vssd1 vccd1 vccd1 _08593_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07544_ _12994_/Q _07531_/A _07568_/A _07532_/A _07538_/X vssd1 vssd1 vccd1 vccd1
+ _12994_/D sky130_fd_sc_hd__o221a_1
XPHY_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07475_ _07475_/A vssd1 vssd1 vccd1 vccd1 _07475_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ _12475_/Q _09207_/X _07536_/X _09208_/X vssd1 vssd1 vccd1 vccd1 _12475_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06426_ _13254_/Q vssd1 vssd1 vccd1 vccd1 _06427_/A sky130_fd_sc_hd__inv_2
XFILLER_50_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09145_ _12506_/Q _09145_/B vssd1 vssd1 vccd1 vccd1 _09146_/B sky130_fd_sc_hd__or2_1
XFILLER_33_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06357_ _12945_/Q vssd1 vssd1 vccd1 vccd1 _06396_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06288_ _06313_/A vssd1 vssd1 vccd1 vccd1 _06288_/X sky130_fd_sc_hd__clkbuf_1
X_09076_ _09180_/C _09180_/D _09179_/A _09179_/B vssd1 vssd1 vccd1 vccd1 _09076_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_136_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08027_ _12876_/Q _08024_/X _07975_/X _08026_/X vssd1 vssd1 vccd1 vccd1 _12876_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_89_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _13152_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09978_ _09981_/A _09978_/B vssd1 vssd1 vccd1 vccd1 _10140_/A sky130_fd_sc_hd__or2_4
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_18_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12489_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08929_ _08929_/A _08929_/B vssd1 vssd1 vccd1 vccd1 _10643_/A sky130_fd_sc_hd__or2_1
XFILLER_58_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11940_ _09648_/Y _12801_/Q _11958_/S vssd1 vssd1 vccd1 vccd1 _11940_/X sky130_fd_sc_hd__mux2_2
XFILLER_18_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11871_ _10210_/Y _12812_/Q _11878_/S vssd1 vssd1 vccd1 vccd1 _11871_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10822_ _12514_/Q _12326_/Q _12515_/Q _12327_/Q vssd1 vssd1 vccd1 vccd1 _10822_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10753_ _10742_/X _10750_/X _06368_/X _10751_/X _10752_/X vssd1 vssd1 vccd1 vccd1
+ _10753_/X sky130_fd_sc_hd__a221o_1
XFILLER_197_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10684_ _12448_/Q _08953_/B _12448_/Q _08953_/B vssd1 vssd1 vccd1 vccd1 _10684_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_199_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12423_ _12620_/CLK _12423_/D vssd1 vssd1 vccd1 vccd1 _12423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12354_ _12570_/CLK _12354_/D vssd1 vssd1 vccd1 vccd1 _12354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ vssd1 vssd1 vccd1 vccd1 _11305_/HI _11305_/LO sky130_fd_sc_hd__conb_1
X_12285_ _12296_/CLK _12285_/D vssd1 vssd1 vccd1 vccd1 _12285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11236_ vssd1 vssd1 vccd1 vccd1 _11236_/HI _11236_/LO sky130_fd_sc_hd__conb_1
XFILLER_136_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11167_ vssd1 vssd1 vccd1 vccd1 _11167_/HI _11167_/LO sky130_fd_sc_hd__conb_1
XFILLER_95_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10118_ _10116_/Y _10018_/X _10117_/Y _10020_/X vssd1 vssd1 vccd1 vccd1 _10128_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_96_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11098_ _11041_/X _11077_/X _06392_/X _11086_/X _11087_/X vssd1 vssd1 vccd1 vccd1
+ _11098_/X sky130_fd_sc_hd__a221o_1
Xinput360 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 input360/X sky130_fd_sc_hd__buf_2
XFILLER_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10049_ _10276_/A vssd1 vssd1 vccd1 vccd1 _10049_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07260_ _07266_/A vssd1 vssd1 vccd1 vccd1 _07260_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_176_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06211_ _06038_/Y _06039_/Y _06046_/B _06210_/X vssd1 vssd1 vccd1 vccd1 _06211_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_192_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07191_ _11516_/X _07160_/A _13115_/Q _07161_/A vssd1 vssd1 vccd1 vccd1 _13115_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06142_ _12736_/Q _12704_/Q _06141_/X vssd1 vssd1 vccd1 vccd1 _06142_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06073_ _12699_/Q vssd1 vssd1 vccd1 vccd1 _06073_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ _12880_/Q _09910_/B vssd1 vssd1 vccd1 vccd1 _09901_/X sky130_fd_sc_hd__or2_1
XFILLER_99_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09832_ _09847_/A _09832_/B vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__or2_1
XFILLER_99_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09763_ _09743_/A _09762_/A _09743_/Y _09762_/Y vssd1 vssd1 vccd1 vccd1 _09769_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06975_ _07026_/A vssd1 vssd1 vccd1 vccd1 _07006_/A sky130_fd_sc_hd__clkbuf_2
X_08714_ _08714_/A vssd1 vssd1 vccd1 vccd1 _08714_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09694_ _09694_/A vssd1 vssd1 vccd1 vccd1 _09694_/Y sky130_fd_sc_hd__inv_2
XPHY_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _08653_/A vssd1 vssd1 vccd1 vccd1 _08645_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08576_ _08715_/A vssd1 vssd1 vccd1 vccd1 _08716_/A sky130_fd_sc_hd__inv_2
XFILLER_82_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07527_ _10527_/B vssd1 vssd1 vccd1 vccd1 _09435_/B sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_136_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12653_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07458_ _07458_/A vssd1 vssd1 vccd1 vccd1 _07458_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06409_ _06412_/A vssd1 vssd1 vccd1 vccd1 _06409_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07389_ _07391_/A vssd1 vssd1 vccd1 vccd1 _07389_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09128_ _12514_/Q _09123_/X _07560_/X _09124_/X vssd1 vssd1 vccd1 vccd1 _12514_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_198_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09059_ _10244_/A vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__buf_6
XFILLER_123_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12070_ _12069_/X _12445_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _12070_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11021_ _12360_/Q _11021_/B vssd1 vssd1 vccd1 vccd1 _11024_/B sky130_fd_sc_hd__nand2_8
XFILLER_132_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12972_ _12974_/CLK _12972_/D vssd1 vssd1 vccd1 vccd1 _12972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11923_ _10274_/Y _12800_/Q _12159_/S vssd1 vssd1 vccd1 vccd1 _11923_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11854_ _11047_/X _11043_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _11854_/X sky130_fd_sc_hd__mux2_1
XPHY_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _12512_/Q _12324_/Q _10804_/Y vssd1 vssd1 vccd1 vccd1 _10807_/A sky130_fd_sc_hd__a21oi_2
XFILLER_198_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11785_ _12120_/X _11784_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11785_/X sky130_fd_sc_hd__mux2_1
XPHY_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10736_ _10736_/A vssd1 vssd1 vccd1 vccd1 _10736_/X sky130_fd_sc_hd__buf_2
XFILLER_14_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ _12429_/Q _12430_/Q vssd1 vssd1 vccd1 vccd1 _10667_/X sky130_fd_sc_hd__and2_1
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12406_ _12410_/CLK _12406_/D vssd1 vssd1 vccd1 vccd1 _12406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10598_ _10607_/A _10598_/B vssd1 vssd1 vccd1 vccd1 _10598_/Y sky130_fd_sc_hd__nor2_1
X_12337_ _12337_/CLK _12337_/D vssd1 vssd1 vccd1 vccd1 _12337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12268_ _10074_/Y _12894_/Q _11857_/X _11858_/X _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12284_/D sky130_fd_sc_hd__mux4_2
X_11219_ vssd1 vssd1 vccd1 vccd1 _11219_/HI _11219_/LO sky130_fd_sc_hd__conb_1
XFILLER_110_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12199_ _10780_/X _11130_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _12199_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06760_ _06758_/X _06759_/X _06758_/X _06759_/X vssd1 vssd1 vccd1 vccd1 _06760_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput190 la_oenb[120] vssd1 vssd1 vccd1 vccd1 input190/X sky130_fd_sc_hd__buf_1
XFILLER_110_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06691_ _11988_/X _11985_/X _11988_/X _11985_/X vssd1 vssd1 vccd1 vccd1 _06691_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08430_ _12776_/Q _08417_/X _07560_/X _08418_/X vssd1 vssd1 vccd1 vccd1 _12776_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08361_ _12803_/Q _08358_/X _07975_/X _08360_/X vssd1 vssd1 vccd1 vccd1 _12803_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07312_ _09184_/A vssd1 vssd1 vccd1 vccd1 _07568_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08292_ _10475_/A _11605_/X _08292_/S vssd1 vssd1 vccd1 vccd1 _12830_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07243_ _07251_/A vssd1 vssd1 vccd1 vccd1 _07243_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07174_ _11523_/X _07160_/X _13122_/Q _07161_/X vssd1 vssd1 vccd1 vccd1 _13122_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06125_ _06125_/A _06125_/B _06125_/C vssd1 vssd1 vccd1 vccd1 _06175_/A sky130_fd_sc_hd__or3_4
XFILLER_132_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06056_ _06056_/A _06241_/A vssd1 vssd1 vccd1 vccd1 _06172_/A sky130_fd_sc_hd__nand2_1
XFILLER_160_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09815_ _09815_/A vssd1 vssd1 vccd1 vccd1 _09823_/B sky130_fd_sc_hd__inv_2
XFILLER_87_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09746_ _09745_/A _09745_/B _09745_/Y vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__a21oi_4
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06958_ _11408_/X _11394_/X vssd1 vssd1 vccd1 vccd1 _06961_/A sky130_fd_sc_hd__or2_1
XFILLER_100_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09677_ _09713_/A _09748_/C vssd1 vssd1 vccd1 vccd1 _09677_/X sky130_fd_sc_hd__or2_1
XFILLER_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06889_ _06916_/A vssd1 vssd1 vccd1 vccd1 _06889_/X sky130_fd_sc_hd__clkbuf_1
XPHY_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _08638_/A vssd1 vssd1 vccd1 vccd1 _08628_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_188_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08559_ _08559_/A vssd1 vssd1 vccd1 vccd1 _12751_/D sky130_fd_sc_hd__inv_2
XPHY_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ _12827_/Q _09179_/C _11578_/S vssd1 vssd1 vccd1 vccd1 _11570_/X sky130_fd_sc_hd__mux2_1
XPHY_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10521_ _10521_/A _10562_/A _10561_/A _10521_/D vssd1 vssd1 vccd1 vccd1 _10526_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_11_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _13241_/CLK _13240_/D _06406_/X vssd1 vssd1 vccd1 vccd1 _13240_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_136_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10452_ _10458_/A _10452_/B _10452_/C vssd1 vssd1 vccd1 vccd1 _10452_/Y sky130_fd_sc_hd__nor3_1
XFILLER_108_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13171_ _13177_/CLK _13171_/D _07011_/X vssd1 vssd1 vccd1 vccd1 _13171_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10383_ _10387_/A _10385_/C _10383_/C vssd1 vssd1 vccd1 vccd1 _10383_/Y sky130_fd_sc_hd__nor3_2
XFILLER_109_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12122_ _12121_/X _12434_/Q _12140_/S vssd1 vssd1 vccd1 vccd1 _12122_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12472_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12053_ _11052_/X _11046_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _12053_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11004_ _11014_/A _11014_/D vssd1 vssd1 vccd1 vccd1 _11004_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12955_ _12955_/CLK _12955_/D vssd1 vssd1 vccd1 vccd1 _12955_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11906_ _08930_/A _10647_/Y _12321_/Q vssd1 vssd1 vccd1 vccd1 _11906_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12886_ _12886_/CLK _12886_/D _07995_/X vssd1 vssd1 vccd1 vccd1 _12886_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ _09945_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11837_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11768_ _09185_/A _11767_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11768_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10719_ _13242_/Q _10738_/A _10699_/A _10737_/A _06430_/X vssd1 vssd1 vccd1 vccd1
+ _10719_/X sky130_fd_sc_hd__o221a_1
XPHY_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11699_ _11396_/X _09180_/C _11703_/S vssd1 vssd1 vccd1 vccd1 _11699_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07930_ _12908_/Q _11497_/X _07932_/S vssd1 vssd1 vccd1 vccd1 _12908_/D sky130_fd_sc_hd__mux2_1
XFILLER_69_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07861_ _07850_/Y _10318_/A _13034_/Q _07824_/Y vssd1 vssd1 vccd1 vccd1 _07866_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_110_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09600_ _09600_/A vssd1 vssd1 vccd1 vccd1 _09600_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06812_ _12022_/X _06789_/X _12022_/X _06789_/X vssd1 vssd1 vccd1 vccd1 _06813_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ _07933_/A vssd1 vssd1 vccd1 vccd1 _07903_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09531_ _09530_/A _09530_/B _09701_/A vssd1 vssd1 vccd1 vccd1 _09531_/Y sky130_fd_sc_hd__o21ai_1
X_06743_ _11991_/X _06691_/X _11991_/X _06691_/X vssd1 vssd1 vccd1 vccd1 _06748_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09462_ _12983_/Q _09436_/X _13006_/Q _09442_/X _09461_/X vssd1 vssd1 vccd1 vccd1
+ _09462_/X sky130_fd_sc_hd__a221o_1
XFILLER_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06674_ _06672_/Y _12051_/X _06673_/X vssd1 vssd1 vccd1 vccd1 _06680_/A sky130_fd_sc_hd__a21oi_2
XFILLER_58_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08413_ _12783_/Q _08401_/X _07990_/X _08403_/X vssd1 vssd1 vccd1 vccd1 _12783_/D
+ sky130_fd_sc_hd__a22o_1
X_09393_ _12395_/D vssd1 vssd1 vccd1 vccd1 _09394_/A sky130_fd_sc_hd__inv_2
XFILLER_33_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08344_ _08352_/A vssd1 vssd1 vccd1 vccd1 _08344_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08275_ _08275_/A vssd1 vssd1 vccd1 vccd1 _08275_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07226_ _07236_/A vssd1 vssd1 vccd1 vccd1 _07226_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07157_ _07167_/A vssd1 vssd1 vccd1 vccd1 _07157_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_105_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06108_ _06108_/A _06108_/B vssd1 vssd1 vccd1 vccd1 _06174_/A sky130_fd_sc_hd__or2_2
X_07088_ _07409_/A vssd1 vssd1 vccd1 vccd1 _08271_/A sky130_fd_sc_hd__buf_4
Xoutput450 _11319_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__clkbuf_2
XFILLER_156_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput461 _11329_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__clkbuf_2
X_06039_ _12711_/Q vssd1 vssd1 vccd1 vccd1 _06039_/Y sky130_fd_sc_hd__inv_2
Xoutput472 _11339_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__clkbuf_2
Xoutput483 _11234_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__clkbuf_2
Xoutput494 _11244_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ _09729_/A vssd1 vssd1 vccd1 vccd1 _09729_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_151_wb_clk_i clkbuf_4_9_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13260_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ _12743_/CLK _12740_/D _08600_/X vssd1 vssd1 vccd1 vccd1 _12740_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12685_/CLK _12671_/D _08789_/X vssd1 vssd1 vccd1 vccd1 _12671_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _10492_/X _12989_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11622_/X sky130_fd_sc_hd__mux2_1
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ _12810_/Q input357/X _11558_/S vssd1 vssd1 vccd1 vccd1 _11553_/X sky130_fd_sc_hd__mux2_1
XPHY_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10504_ _12509_/Q _09147_/X _12509_/Q _09147_/X vssd1 vssd1 vccd1 vccd1 _10504_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_13_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11484_ _10325_/Y _09185_/C _11487_/S vssd1 vssd1 vccd1 vccd1 _11484_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13223_ _13223_/CLK _13223_/D _06554_/X vssd1 vssd1 vccd1 vccd1 _13223_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10435_ _10433_/B _10433_/C _10433_/A vssd1 vssd1 vccd1 vccd1 _10436_/C sky130_fd_sc_hd__o21a_1
XFILLER_100_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13154_ _13154_/CLK _13154_/D _07063_/X vssd1 vssd1 vccd1 vccd1 _13154_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_100_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10366_ _10367_/B _10363_/A _12911_/Q _10365_/B _10350_/X vssd1 vssd1 vccd1 vccd1
+ _10366_/X sky130_fd_sc_hd__o221a_1
XFILLER_152_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12105_ _12431_/Q _10668_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12105_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13085_ _12167_/X _13085_/D _07274_/X vssd1 vssd1 vccd1 vccd1 _13085_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10297_ _10295_/Y _10032_/X _10296_/Y _10028_/X vssd1 vssd1 vccd1 vccd1 _10297_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_151_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12036_ _11070_/X _11065_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12938_ _12939_/CLK _12938_/D vssd1 vssd1 vccd1 vccd1 _12938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _12886_/CLK _12869_/D _08043_/X vssd1 vssd1 vccd1 vccd1 _12869_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06390_ _06382_/X _12216_/X _06375_/X _06389_/X vssd1 vssd1 vccd1 vccd1 _13245_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08060_ _12862_/Q _08040_/A _07309_/X _08041_/A vssd1 vssd1 vccd1 vccd1 _12862_/D
+ sky130_fd_sc_hd__a22o_1
X_07011_ _07024_/A vssd1 vssd1 vccd1 vccd1 _07011_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08962_ _08962_/A vssd1 vssd1 vccd1 vccd1 _08962_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07913_ _07917_/A vssd1 vssd1 vccd1 vccd1 _07913_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08893_ _12612_/Q vssd1 vssd1 vccd1 vccd1 _08893_/X sky130_fd_sc_hd__buf_2
XFILLER_190_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07844_ _13031_/Q _10380_/B _12836_/Q vssd1 vssd1 vccd1 vccd1 _07867_/A sky130_fd_sc_hd__o21ai_1
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07775_ _07775_/A vssd1 vssd1 vccd1 vccd1 _07775_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09514_ _09514_/A vssd1 vssd1 vccd1 vccd1 _09514_/Y sky130_fd_sc_hd__inv_2
X_06726_ _12033_/X _06724_/B _06724_/X vssd1 vssd1 vccd1 vccd1 _06726_/X sky130_fd_sc_hd__a21bo_1
XFILLER_197_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09445_ _12966_/Q _09440_/X _13002_/Q _09442_/X _09444_/X vssd1 vssd1 vccd1 vccd1
+ _09445_/X sky130_fd_sc_hd__a221o_1
X_06657_ _06690_/A vssd1 vssd1 vccd1 vccd1 _06657_/X sky130_fd_sc_hd__clkbuf_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ _12407_/Q vssd1 vssd1 vccd1 vccd1 _09376_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06588_ _12202_/X _12201_/X _06587_/X vssd1 vssd1 vccd1 vccd1 _06588_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08327_ _08372_/A vssd1 vssd1 vccd1 vccd1 _08339_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08258_ _12840_/Q _08251_/X _07296_/X _11417_/S vssd1 vssd1 vccd1 vccd1 _12840_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07209_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07209_/X sky130_fd_sc_hd__clkbuf_1
X_08189_ _13114_/Q _08176_/Y _13134_/Q _10460_/A _08188_/X vssd1 vssd1 vccd1 vccd1
+ _08190_/D sky130_fd_sc_hd__o221a_1
XFILLER_106_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10220_ _12631_/Q vssd1 vssd1 vccd1 vccd1 _10220_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10151_ _10151_/A vssd1 vssd1 vccd1 vccd1 _10151_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10082_ _10081_/Y _10137_/A _09896_/Y _10003_/A vssd1 vssd1 vccd1 vccd1 _10088_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10984_ _12538_/Q _12350_/Q _10975_/Y _10980_/Y vssd1 vssd1 vccd1 vccd1 _10985_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12723_ _13162_/CLK _12723_/D _08645_/X vssd1 vssd1 vccd1 vccd1 _12723_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ _13264_/CLK _12654_/D _08834_/X vssd1 vssd1 vccd1 vccd1 _12654_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _10476_/X _10794_/D _11610_/S vssd1 vssd1 vccd1 vccd1 _11605_/X sky130_fd_sc_hd__mux2_1
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _12586_/CLK _12585_/D vssd1 vssd1 vccd1 vccd1 _12585_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11536_ _12825_/Q _09180_/A _11543_/S vssd1 vssd1 vccd1 vccd1 _11536_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11467_ _12910_/Q _09179_/A _11469_/S vssd1 vssd1 vccd1 vccd1 _11467_/X sky130_fd_sc_hd__mux2_1
X_13206_ _13208_/CLK _13206_/D _06718_/X vssd1 vssd1 vccd1 vccd1 _13206_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10418_ _10418_/A _10418_/B vssd1 vssd1 vccd1 vccd1 _10420_/B sky130_fd_sc_hd__or2_2
XFILLER_171_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11398_ _10605_/Y _12409_/D _11404_/S vssd1 vssd1 vccd1 vccd1 _11398_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13137_ _12168_/X _13137_/D _07135_/X vssd1 vssd1 vccd1 vccd1 _13137_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10349_ _10371_/A _10349_/B _10349_/C vssd1 vssd1 vccd1 vccd1 _10349_/Y sky130_fd_sc_hd__nor3_1
XFILLER_135_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13068_ _12165_/X _13068_/D _07335_/X vssd1 vssd1 vccd1 vccd1 _13068_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12019_ _11092_/X _11085_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _12019_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ _09186_/A vssd1 vssd1 vccd1 vccd1 _07560_/X sky130_fd_sc_hd__buf_4
XFILLER_98_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06511_ _12162_/X vssd1 vssd1 vccd1 vccd1 _06511_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07491_ _07933_/A vssd1 vssd1 vccd1 vccd1 _07749_/A sky130_fd_sc_hd__buf_6
XFILLER_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09230_ _09247_/A _11675_/S vssd1 vssd1 vccd1 vccd1 _09232_/A sky130_fd_sc_hd__nand2_1
X_06442_ _11900_/X vssd1 vssd1 vccd1 vccd1 _06444_/A sky130_fd_sc_hd__inv_2
XFILLER_167_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09161_ _11630_/X _09154_/X _12505_/Q _09156_/X vssd1 vssd1 vccd1 vccd1 _12505_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06373_ _06416_/A vssd1 vssd1 vccd1 vccd1 _06391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08112_ _13117_/Q vssd1 vssd1 vccd1 vccd1 _08112_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09092_ _09116_/A vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08043_ _08051_/A vssd1 vssd1 vccd1 vccd1 _08043_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09994_ _08790_/Y _09993_/X _06258_/Y _09972_/X _09991_/X vssd1 vssd1 vccd1 vccd1
+ _09994_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08945_ _12445_/Q _12446_/Q vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__or2_1
XFILLER_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08876_ _12612_/Q vssd1 vssd1 vccd1 vccd1 _08898_/A sky130_fd_sc_hd__inv_2
XFILLER_56_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07827_ _13026_/Q vssd1 vssd1 vccd1 vccd1 _07827_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07758_ _12584_/Q _07758_/B vssd1 vssd1 vccd1 vccd1 _07759_/B sky130_fd_sc_hd__or2_1
XFILLER_72_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06709_ _06750_/A vssd1 vssd1 vccd1 vccd1 _06709_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_197_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07689_ _07668_/B _07689_/B _07689_/C _07689_/D vssd1 vssd1 vccd1 vccd1 _07690_/B
+ sky130_fd_sc_hd__and4b_1
X_09428_ _12415_/D vssd1 vssd1 vccd1 vccd1 _09428_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09359_ _09354_/Y _12400_/Q _09355_/Y _12415_/Q _09358_/X vssd1 vssd1 vccd1 vccd1
+ _09359_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12370_ _12376_/CLK _12370_/D vssd1 vssd1 vccd1 vccd1 _12370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11321_ vssd1 vssd1 vccd1 vccd1 _11321_/HI _11321_/LO sky130_fd_sc_hd__conb_1
XFILLER_193_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11252_ vssd1 vssd1 vccd1 vccd1 _11252_/HI _11252_/LO sky130_fd_sc_hd__conb_1
XFILLER_107_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10203_ _09569_/Y _10166_/X _10202_/Y _10168_/X vssd1 vssd1 vccd1 vccd1 _10203_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11183_ vssd1 vssd1 vccd1 vccd1 _11183_/HI _11183_/LO sky130_fd_sc_hd__conb_1
XFILLER_106_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10134_ _10134_/A vssd1 vssd1 vccd1 vccd1 _10134_/X sky130_fd_sc_hd__buf_2
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10065_ _12773_/Q vssd1 vssd1 vccd1 vccd1 _10065_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10967_ _10977_/A _10977_/B _10977_/D _10966_/Y vssd1 vssd1 vccd1 vccd1 _10967_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_189_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12706_ _12707_/CLK _12706_/D _08689_/X vssd1 vssd1 vccd1 vccd1 _12706_/Q sky130_fd_sc_hd__dfrtp_2
X_10898_ _12527_/Q vssd1 vssd1 vccd1 vccd1 _10900_/A sky130_fd_sc_hd__inv_2
XFILLER_188_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ _13162_/CLK _12637_/D _08875_/X vssd1 vssd1 vccd1 vccd1 _12637_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12568_ _12570_/CLK _12568_/D vssd1 vssd1 vccd1 vccd1 _12568_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11519_ _12808_/Q _09186_/A _11522_/S vssd1 vssd1 vccd1 vccd1 _11519_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12499_ _12586_/CLK _12499_/D vssd1 vssd1 vccd1 vccd1 _12499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06991_ _06995_/A _06995_/B vssd1 vssd1 vccd1 vccd1 _06991_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08730_ _11823_/X _08592_/A _12689_/Q _08593_/A vssd1 vssd1 vccd1 vccd1 _12689_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08661_ _08669_/A vssd1 vssd1 vccd1 vccd1 _08661_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07612_ _11618_/X _07610_/X _12973_/Q _07611_/X _07583_/X vssd1 vssd1 vccd1 vccd1
+ _12973_/D sky130_fd_sc_hd__o221a_1
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08592_ _08592_/A vssd1 vssd1 vccd1 vccd1 _08592_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07543_ _12995_/Q _07531_/A _09226_/B _07532_/A _07538_/X vssd1 vssd1 vccd1 vccd1
+ _12995_/D sky130_fd_sc_hd__o221a_1
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07474_ _07474_/A vssd1 vssd1 vccd1 vccd1 _07474_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09213_ _12476_/Q _09207_/X _07545_/X _09208_/X vssd1 vssd1 vccd1 vccd1 _12476_/D
+ sky130_fd_sc_hd__a22o_1
X_06425_ _06425_/A vssd1 vssd1 vccd1 vccd1 _10738_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09144_ _12505_/Q _09144_/B vssd1 vssd1 vccd1 vccd1 _09145_/B sky130_fd_sc_hd__or2_1
X_06356_ _13254_/Q vssd1 vssd1 vccd1 vccd1 _06356_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_33_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09075_ _09083_/A vssd1 vssd1 vccd1 vccd1 _09247_/A sky130_fd_sc_hd__inv_2
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06287_ _06416_/A vssd1 vssd1 vccd1 vccd1 _06313_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08026_ _08041_/A vssd1 vssd1 vccd1 vccd1 _08026_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09977_ _12787_/Q vssd1 vssd1 vccd1 vccd1 _09977_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08928_ _08928_/A _10636_/A vssd1 vssd1 vccd1 vccd1 _08929_/B sky130_fd_sc_hd__or2_1
XFILLER_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08859_ _08849_/X _06316_/X _08852_/X _12645_/Q vssd1 vssd1 vccd1 vccd1 _12645_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_55_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_58_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12992_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11870_ _10190_/Y _12320_/Q _12312_/Q vssd1 vssd1 vccd1 vccd1 _11870_/X sky130_fd_sc_hd__mux2_2
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10821_ _10821_/A _10821_/B _10821_/C vssd1 vssd1 vccd1 vccd1 _10828_/A sky130_fd_sc_hd__nor3_4
XFILLER_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10752_ _12089_/X vssd1 vssd1 vccd1 vccd1 _10752_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10683_ _12447_/Q _08946_/B _08953_/B vssd1 vssd1 vccd1 vccd1 _10683_/X sky130_fd_sc_hd__a21bo_1
XFILLER_197_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12422_ _12422_/CLK _12422_/D vssd1 vssd1 vccd1 vccd1 _12422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12353_ _12353_/CLK _12353_/D vssd1 vssd1 vccd1 vccd1 _12353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11304_ vssd1 vssd1 vccd1 vccd1 _11304_/HI _11304_/LO sky130_fd_sc_hd__conb_1
X_12284_ _12284_/CLK _12284_/D vssd1 vssd1 vccd1 vccd1 _12284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11235_ vssd1 vssd1 vccd1 vccd1 _11235_/HI _11235_/LO sky130_fd_sc_hd__conb_1
XFILLER_107_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11166_ vssd1 vssd1 vccd1 vccd1 _11166_/HI _11166_/LO sky130_fd_sc_hd__conb_1
XFILLER_136_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10117_ _12881_/Q vssd1 vssd1 vccd1 vccd1 _10117_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13235_/CLK
+ sky130_fd_sc_hd__clkbuf_1
X_11097_ _10773_/X _11075_/X _13246_/Q _11083_/X _11084_/X vssd1 vssd1 vccd1 vccd1
+ _11097_/X sky130_fd_sc_hd__a221o_1
XFILLER_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput350 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 _10794_/A sky130_fd_sc_hd__buf_4
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput361 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _09293_/A sky130_fd_sc_hd__buf_1
X_10048_ _10151_/A vssd1 vssd1 vccd1 vccd1 _10276_/A sky130_fd_sc_hd__inv_2
XFILLER_76_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _11104_/X _11096_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _11999_/X sky130_fd_sc_hd__mux2_2
XFILLER_44_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06210_ _06209_/A _06209_/B _06183_/X _06170_/X _06209_/X vssd1 vssd1 vccd1 vccd1
+ _06210_/X sky130_fd_sc_hd__o311a_1
XFILLER_192_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07190_ _07206_/A vssd1 vssd1 vccd1 vccd1 _07190_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_129_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06141_ _12736_/Q _12704_/Q _12735_/Q _12703_/Q vssd1 vssd1 vccd1 vccd1 _06141_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06072_ _12731_/Q vssd1 vssd1 vccd1 vccd1 _06072_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09900_ _12657_/Q vssd1 vssd1 vccd1 vccd1 _09900_/Y sky130_fd_sc_hd__inv_2
X_09831_ _09847_/A _09832_/B vssd1 vssd1 vccd1 vccd1 _09831_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09762_ _09762_/A vssd1 vssd1 vccd1 vccd1 _09762_/Y sky130_fd_sc_hd__inv_2
X_06974_ _06886_/X _12187_/X _06887_/X _13178_/Q vssd1 vssd1 vccd1 vccd1 _13178_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08713_ _11830_/X _08700_/X _12696_/Q _08701_/X vssd1 vssd1 vccd1 vccd1 _12696_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09693_ _09686_/X _09692_/X _09686_/X _09692_/X vssd1 vssd1 vccd1 vccd1 _09694_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08644_ _11933_/X _08639_/X _12724_/Q _08640_/X vssd1 vssd1 vccd1 vccd1 _12724_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08575_ _08592_/A vssd1 vssd1 vccd1 vccd1 _08575_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07526_ _13001_/Q vssd1 vssd1 vccd1 vccd1 _09019_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_81_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07457_ _11464_/X _07444_/X _13023_/Q _07445_/X vssd1 vssd1 vccd1 vccd1 _13023_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06408_ _06403_/X _12206_/X _06396_/X _06407_/X vssd1 vssd1 vccd1 vccd1 _13240_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07388_ _11424_/X _07384_/X _13048_/Q _07385_/X vssd1 vssd1 vccd1 vccd1 _13048_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09127_ _12515_/Q _09123_/X _07558_/X _09124_/X vssd1 vssd1 vccd1 vccd1 _12515_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06339_ _06115_/Y _06116_/Y _12720_/Q _12688_/Q vssd1 vssd1 vccd1 vccd1 _06339_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09058_ _09058_/A _12148_/X vssd1 vssd1 vccd1 vccd1 _12559_/D sky130_fd_sc_hd__nor2b_1
XFILLER_68_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08009_ _12882_/Q _07996_/X _07293_/X _07998_/X vssd1 vssd1 vccd1 vccd1 _12882_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11020_ _11021_/B _11020_/B vssd1 vssd1 vccd1 vccd1 _12359_/D sky130_fd_sc_hd__nor2_1
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12971_ _12974_/CLK _12971_/D vssd1 vssd1 vccd1 vccd1 _12971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11922_ _11921_/X _12442_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _11922_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _11039_/X _11036_/Y _12186_/S vssd1 vssd1 vccd1 vccd1 _11853_/X sky130_fd_sc_hd__mux2_2
XPHY_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10804_ _12512_/Q _12324_/Q vssd1 vssd1 vccd1 vccd1 _10804_/Y sky130_fd_sc_hd__nor2_1
X_11784_ _09244_/B _11783_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11784_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10735_ _13252_/Q vssd1 vssd1 vccd1 vccd1 _10736_/A sky130_fd_sc_hd__inv_2
XFILLER_201_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10666_ _12429_/Q vssd1 vssd1 vccd1 vccd1 _10666_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12405_ _12410_/CLK _12405_/D vssd1 vssd1 vccd1 vccd1 _12405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10597_ _12407_/D _11403_/S _10599_/A _10588_/A vssd1 vssd1 vccd1 vccd1 _10598_/B
+ sky130_fd_sc_hd__o22a_1
X_12336_ _12337_/CLK _12336_/D vssd1 vssd1 vccd1 vccd1 _12336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12267_ _10055_/X _12893_/Q _11855_/X _11856_/X _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12283_/D sky130_fd_sc_hd__mux4_2
XFILLER_142_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11218_ vssd1 vssd1 vccd1 vccd1 _11218_/HI _11218_/LO sky130_fd_sc_hd__conb_1
X_12198_ _10748_/X _10749_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _12198_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11149_ vssd1 vssd1 vccd1 vccd1 _11149_/HI _11149_/LO sky130_fd_sc_hd__conb_1
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput180 la_oenb[111] vssd1 vssd1 vccd1 vccd1 input180/X sky130_fd_sc_hd__buf_1
Xinput191 la_oenb[121] vssd1 vssd1 vccd1 vccd1 input191/X sky130_fd_sc_hd__buf_1
XFILLER_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06690_ _06690_/A vssd1 vssd1 vccd1 vccd1 _06690_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08360_ _08375_/A vssd1 vssd1 vccd1 vccd1 _08360_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07311_ _07330_/A vssd1 vssd1 vccd1 vccd1 _07311_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_3_wb_clk_i _12844_/CLK vssd1 vssd1 vccd1 vccd1 _12169_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_147_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08291_ _08296_/A vssd1 vssd1 vccd1 vccd1 _08291_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07242_ _11563_/X _07233_/X _13098_/Q _07234_/X vssd1 vssd1 vccd1 vccd1 _13098_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07173_ _07183_/A vssd1 vssd1 vccd1 vccd1 _07173_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06124_ _06115_/Y _06116_/Y _06122_/Y _06123_/X vssd1 vssd1 vccd1 vccd1 _06125_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06055_ _06053_/Y _06054_/Y _12737_/Q _12705_/Q vssd1 vssd1 vccd1 vccd1 _06241_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_114_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09814_ _09826_/A _09813_/X _09826_/A _09813_/X vssd1 vssd1 vccd1 vccd1 _09815_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ _09745_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09745_/Y sky130_fd_sc_hd__nor2_4
X_06957_ _13179_/Q vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__inv_2
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09676_ _09632_/B _09714_/A _09611_/B _09674_/Y _09675_/X vssd1 vssd1 vccd1 vccd1
+ _09748_/C sky130_fd_sc_hd__o311a_1
X_06888_ _06886_/X _12188_/X _06887_/X _13188_/Q vssd1 vssd1 vccd1 vccd1 _13188_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _08642_/A vssd1 vssd1 vccd1 vccd1 _08638_/A sky130_fd_sc_hd__clkbuf_2
XPHY_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _08552_/X _08553_/Y _08558_/S vssd1 vssd1 vccd1 vccd1 _08559_/A sky130_fd_sc_hd__mux2_1
XPHY_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07509_ _09228_/B _07497_/Y _07522_/B _11982_/X _07508_/Y vssd1 vssd1 vccd1 vccd1
+ _07510_/B sky130_fd_sc_hd__o32a_1
XPHY_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08489_ _08453_/Y _07815_/X _13069_/Q _10390_/A vssd1 vssd1 vccd1 vccd1 _08489_/X
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ _10579_/A _12402_/D _10520_/C _12400_/D vssd1 vssd1 vccd1 vccd1 _10521_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_156_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10451_ _10449_/B _10455_/D _10455_/A vssd1 vssd1 vccd1 vccd1 _10452_/C sky130_fd_sc_hd__o21a_1
XFILLER_183_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13170_ _13170_/CLK _13170_/D _07014_/X vssd1 vssd1 vccd1 vccd1 _13170_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10382_ _10380_/B _10380_/C _10380_/A vssd1 vssd1 vccd1 vccd1 _10383_/C sky130_fd_sc_hd__o21a_1
XFILLER_151_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12121_ _10671_/X _09313_/X _12121_/S vssd1 vssd1 vccd1 vccd1 _12121_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ _10774_/X _11126_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _12052_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11003_ _10980_/B _11000_/X _10980_/A _11000_/X _11002_/Y vssd1 vssd1 vccd1 vccd1
+ _11014_/D sky130_fd_sc_hd__o221a_2
XFILLER_46_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_wb_clk_i _12960_/CLK vssd1 vssd1 vccd1 vccd1 _12961_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12954_ _12957_/CLK _12954_/D vssd1 vssd1 vccd1 vccd1 _12954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11905_ _08929_/A _10644_/X _12321_/Q vssd1 vssd1 vccd1 vccd1 _11905_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ _12886_/CLK _12885_/D _08000_/X vssd1 vssd1 vccd1 vccd1 _12885_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _09944_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11836_/X sky130_fd_sc_hd__mux2_1
XPHY_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11767_ _12111_/X _12476_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11767_/X sky130_fd_sc_hd__mux2_1
XPHY_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10718_ _13243_/Q _10738_/A _11033_/A _10717_/X _06430_/X vssd1 vssd1 vccd1 vccd1
+ _10781_/A sky130_fd_sc_hd__o221a_1
XPHY_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11698_ _11697_/X _11399_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12391_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10649_ _11906_/X _10649_/B vssd1 vssd1 vccd1 vccd1 _10649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12319_ _12987_/CLK _12319_/D vssd1 vssd1 vccd1 vccd1 _12319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07860_ _12894_/Q vssd1 vssd1 vccd1 vccd1 _10318_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_111_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06811_ _11881_/X _06807_/Y _06810_/Y vssd1 vssd1 vccd1 vccd1 _06813_/A sky130_fd_sc_hd__o21a_1
X_07791_ _07522_/B _07520_/A _07562_/A _07616_/X _07790_/X vssd1 vssd1 vccd1 vccd1
+ _12925_/D sky130_fd_sc_hd__o311a_1
XFILLER_96_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06742_ _06740_/X _06741_/X _06740_/X _06741_/X vssd1 vssd1 vccd1 vccd1 _06748_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_09530_ _09530_/A _09530_/B vssd1 vssd1 vccd1 vccd1 _09530_/X sky130_fd_sc_hd__and2_1
XFILLER_97_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09461_ _12931_/Q _09438_/X _12999_/Q _09451_/X _09460_/X vssd1 vssd1 vccd1 vccd1
+ _09461_/X sky130_fd_sc_hd__a221o_1
XFILLER_97_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06673_ _11897_/X _06643_/X _11897_/X _06643_/X vssd1 vssd1 vccd1 vccd1 _06673_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_184_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08412_ _08420_/A vssd1 vssd1 vccd1 vccd1 _08412_/X sky130_fd_sc_hd__clkbuf_1
X_09392_ _12463_/Q _10520_/C _09375_/Y _12407_/D _09391_/X vssd1 vssd1 vccd1 vccd1
+ _09402_/B sky130_fd_sc_hd__o221a_1
XFILLER_149_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08343_ _12809_/Q _11584_/X _08349_/S vssd1 vssd1 vccd1 vccd1 _12809_/D sky130_fd_sc_hd__mux2_1
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08274_ _08273_/Y input12/X _08273_/Y input12/X vssd1 vssd1 vccd1 vccd1 _08274_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_165_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07225_ _11570_/X _07218_/X _13105_/Q _07219_/X vssd1 vssd1 vccd1 vccd1 _13105_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07156_ _11530_/X _07145_/X _13129_/Q _07146_/X vssd1 vssd1 vccd1 vccd1 _13129_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06107_ _12723_/Q _12691_/Q _06105_/Y _06106_/Y vssd1 vssd1 vccd1 vccd1 _06108_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07087_ _10527_/A _07515_/A _09434_/B _09073_/A vssd1 vssd1 vccd1 vccd1 _07409_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput440 _12844_/Q vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput451 _11320_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__clkbuf_2
X_06038_ _12743_/Q vssd1 vssd1 vccd1 vccd1 _06038_/Y sky130_fd_sc_hd__inv_2
Xoutput462 _11330_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__clkbuf_2
Xoutput473 _11340_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__clkbuf_2
Xoutput484 _11235_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput495 _11245_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07989_ _08004_/A vssd1 vssd1 vccd1 vccd1 _07989_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09728_ _09721_/Y _09727_/X _09721_/Y _09727_/X vssd1 vssd1 vccd1 vccd1 _09729_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09659_ _09659_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _09659_/X sky130_fd_sc_hd__or2_1
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12682_/CLK _12670_/D _08793_/X vssd1 vssd1 vccd1 vccd1 _12670_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11621_ _10491_/X _12988_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11621_/X sky130_fd_sc_hd__mux2_1
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_120_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 _12685_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ _12809_/Q _09185_/B _11558_/S vssd1 vssd1 vccd1 vccd1 _11552_/X sky130_fd_sc_hd__mux2_1
XPHY_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10503_ _12508_/Q _09147_/B _09147_/X vssd1 vssd1 vccd1 vccd1 _10503_/X sky130_fd_sc_hd__a21bo_1
XFILLER_52_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11483_ _10321_/X _09185_/D _11487_/S vssd1 vssd1 vccd1 vccd1 _11483_/X sky130_fd_sc_hd__mux2_1
XPHY_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13222_ _13236_/CLK _13222_/D _06560_/X vssd1 vssd1 vccd1 vccd1 _13222_/Q sky130_fd_sc_hd__dfrtp_1
X_10434_ _10439_/C vssd1 vssd1 vccd1 vccd1 _10436_/B sky130_fd_sc_hd__inv_2
XFILLER_100_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10365_ _10371_/A _10365_/B _10365_/C vssd1 vssd1 vccd1 vccd1 _10365_/Y sky130_fd_sc_hd__nor3_1
XFILLER_83_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13153_ _13154_/CLK _13153_/D _07066_/X vssd1 vssd1 vccd1 vccd1 _13153_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12104_ _12103_/X _12430_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12104_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13084_ _12167_/X _13084_/D _07276_/X vssd1 vssd1 vccd1 vccd1 _13084_/Q sky130_fd_sc_hd__dfrtp_4
X_10296_ _12859_/Q vssd1 vssd1 vccd1 vccd1 _10296_/Y sky130_fd_sc_hd__inv_2
X_12035_ _11116_/X _11104_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _12035_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12937_ _12937_/CLK _12937_/D vssd1 vssd1 vccd1 vccd1 _12937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _12868_/CLK _12868_/D _08045_/X vssd1 vssd1 vccd1 vccd1 _12868_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11819_ _11818_/X _12096_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12448_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12799_ _12801_/CLK _12799_/D _08368_/X vssd1 vssd1 vccd1 vccd1 _12799_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_193_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07010_ _07026_/A vssd1 vssd1 vccd1 vccd1 _07024_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_161_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08961_ _08962_/A vssd1 vssd1 vccd1 vccd1 _08961_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07912_ _12916_/Q _11505_/X _07918_/S vssd1 vssd1 vccd1 vccd1 _12916_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08892_ _08897_/A vssd1 vssd1 vccd1 vccd1 _08892_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07843_ _12915_/Q vssd1 vssd1 vccd1 vccd1 _10380_/B sky130_fd_sc_hd__inv_2
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07774_ _12934_/Q _07768_/A _12935_/Q _07769_/X _07569_/X vssd1 vssd1 vccd1 vccd1
+ _12935_/D sky130_fd_sc_hd__a221o_1
X_09513_ _13172_/Q _13171_/Q _09526_/A _09526_/B vssd1 vssd1 vccd1 vccd1 _09514_/A
+ sky130_fd_sc_hd__o22a_1
X_06725_ _12009_/X _12035_/X _06724_/X vssd1 vssd1 vccd1 vccd1 _06725_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06656_ _06766_/A vssd1 vssd1 vccd1 vccd1 _06690_/A sky130_fd_sc_hd__clkbuf_2
X_09444_ _12571_/Q _07519_/B _12994_/Q _09451_/A vssd1 vssd1 vccd1 vccd1 _09444_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09375_ _12455_/Q vssd1 vssd1 vccd1 vccd1 _09375_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06587_ _12200_/X _06587_/B vssd1 vssd1 vccd1 vccd1 _06587_/X sky130_fd_sc_hd__or2_1
XFILLER_178_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08326_ _12816_/Q _11591_/X _08335_/S vssd1 vssd1 vccd1 vccd1 _12816_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08257_ _08257_/A vssd1 vssd1 vccd1 vccd1 _08257_/X sky130_fd_sc_hd__clkbuf_1
X_07208_ _07253_/A vssd1 vssd1 vccd1 vccd1 _07221_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_165_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08188_ _13126_/Q _08187_/X _13126_/Q _08187_/X vssd1 vssd1 vccd1 vccd1 _08188_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07139_ _07154_/A vssd1 vssd1 vccd1 vccd1 _07152_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10150_ _10150_/A _11977_/X vssd1 vssd1 vccd1 vccd1 _10150_/Y sky130_fd_sc_hd__nor2b_1
X_10081_ _12847_/Q vssd1 vssd1 vccd1 vccd1 _10081_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10983_ _11000_/B vssd1 vssd1 vccd1 vccd1 _10983_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12722_ _13162_/CLK _12722_/D _08647_/X vssd1 vssd1 vccd1 vccd1 _12722_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ _12653_/CLK _12653_/D _08836_/X vssd1 vssd1 vccd1 vccd1 _12653_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ _10474_/Y _10792_/A _11610_/S vssd1 vssd1 vccd1 vccd1 _11604_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _12586_/CLK _12584_/D vssd1 vssd1 vccd1 vccd1 _12584_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11535_ _12824_/Q _09180_/B _11543_/S vssd1 vssd1 vccd1 vccd1 _11535_/X sky130_fd_sc_hd__mux2_1
XPHY_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11466_ _12909_/Q _09179_/B _11469_/S vssd1 vssd1 vccd1 vccd1 _11466_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13205_ _13205_/CLK _13205_/D _06722_/X vssd1 vssd1 vccd1 vccd1 _13205_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10417_ _10415_/A _10415_/B _10416_/Y _10411_/A vssd1 vssd1 vccd1 vccd1 _10417_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_174_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11397_ _10606_/X _12410_/D _11403_/S vssd1 vssd1 vccd1 vccd1 _11397_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ _12168_/X _13136_/D _07137_/X vssd1 vssd1 vccd1 vccd1 _13136_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_124_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10348_ _10346_/B _10346_/C _10346_/A vssd1 vssd1 vccd1 vccd1 _10349_/C sky130_fd_sc_hd__o21a_1
XFILLER_152_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13067_ _12165_/X _13067_/D _07337_/X vssd1 vssd1 vccd1 vccd1 _13067_/Q sky130_fd_sc_hd__dfrtp_1
X_10279_ _13021_/Q _10276_/X _13054_/Q _10277_/X vssd1 vssd1 vccd1 vccd1 _10279_/X
+ sky130_fd_sc_hd__a22o_1
X_12018_ _11091_/X _11082_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _12018_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06510_ _11959_/X vssd1 vssd1 vccd1 vccd1 _06510_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07490_ _11451_/X _07459_/A _13010_/Q _07460_/A vssd1 vssd1 vccd1 vccd1 _13010_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06441_ _13235_/Q vssd1 vssd1 vccd1 vccd1 _06441_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09160_ _11631_/X _09154_/X _12506_/Q _09156_/X vssd1 vssd1 vccd1 vccd1 _12506_/D
+ sky130_fd_sc_hd__a22o_1
X_06372_ _06361_/X _12226_/X _06358_/X _06371_/X vssd1 vssd1 vccd1 vccd1 _13250_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08111_ _08105_/Y _12808_/Q _13118_/Q _10415_/A _08110_/X vssd1 vssd1 vccd1 vccd1
+ _08132_/A sky130_fd_sc_hd__a221o_1
XFILLER_30_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09091_ _09124_/A vssd1 vssd1 vccd1 vccd1 _09116_/A sky130_fd_sc_hd__buf_4
XFILLER_147_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08042_ _12870_/Q _08040_/X _07997_/X _08041_/X vssd1 vssd1 vccd1 vccd1 _12870_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09993_ _10003_/A vssd1 vssd1 vccd1 vccd1 _09993_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ _08944_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _09311_/A sky130_fd_sc_hd__nand2_4
XFILLER_85_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08875_ _08882_/A vssd1 vssd1 vccd1 vccd1 _08875_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07826_ _07820_/Y _07821_/X _13009_/Q _07822_/Y _07825_/X vssd1 vssd1 vccd1 vccd1
+ _07842_/A sky130_fd_sc_hd__a221o_1
XFILLER_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07757_ _12583_/Q _07757_/B vssd1 vssd1 vccd1 vccd1 _07758_/B sky130_fd_sc_hd__or2_1
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06708_ _06766_/A vssd1 vssd1 vccd1 vccd1 _06750_/A sky130_fd_sc_hd__clkbuf_2
X_07688_ _07688_/A vssd1 vssd1 vccd1 vccd1 _07688_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09427_ _12466_/Q _09415_/Y _12467_/Q _09426_/X vssd1 vssd1 vccd1 vccd1 _09427_/X
+ sky130_fd_sc_hd__o211a_1
X_06639_ _12198_/X _10765_/A vssd1 vssd1 vccd1 vccd1 _06639_/X sky130_fd_sc_hd__or2_1
XFILLER_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09358_ _12460_/Q _09356_/Y _09357_/Y _12416_/Q vssd1 vssd1 vccd1 vccd1 _09358_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08309_ _08353_/S vssd1 vssd1 vccd1 vccd1 _08321_/S sky130_fd_sc_hd__buf_2
XFILLER_139_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09289_ _07711_/A _09278_/Y _09027_/B _09288_/Y _09262_/X vssd1 vssd1 vccd1 vccd1
+ _12308_/D sky130_fd_sc_hd__o221ai_1
XFILLER_138_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11320_ vssd1 vssd1 vccd1 vccd1 _11320_/HI _11320_/LO sky130_fd_sc_hd__conb_1
XFILLER_181_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11251_ vssd1 vssd1 vccd1 vccd1 _11251_/HI _11251_/LO sky130_fd_sc_hd__conb_1
XFILLER_140_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10202_ _12646_/Q vssd1 vssd1 vccd1 vccd1 _10202_/Y sky130_fd_sc_hd__inv_2
X_11182_ vssd1 vssd1 vccd1 vccd1 _11182_/HI _11182_/LO sky130_fd_sc_hd__conb_1
XFILLER_122_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10133_ _11969_/S _10527_/C _09982_/D _12840_/Q _10132_/X vssd1 vssd1 vccd1 vccd1
+ _10133_/X sky130_fd_sc_hd__a41o_1
XFILLER_192_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10064_ _12862_/Q vssd1 vssd1 vccd1 vccd1 _10064_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10966_ _12535_/Q _12347_/Q _10965_/X vssd1 vssd1 vccd1 vccd1 _10966_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_189_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12705_ _12707_/CLK _12705_/D _08691_/X vssd1 vssd1 vccd1 vccd1 _12705_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10897_ _10895_/A _10921_/A _10895_/Y _10896_/Y vssd1 vssd1 vccd1 vccd1 _12338_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_188_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12636_ _13162_/CLK _12636_/D _08880_/X vssd1 vssd1 vccd1 vccd1 _12636_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12567_ _12570_/CLK _12567_/D vssd1 vssd1 vccd1 vccd1 _12567_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11518_ _12807_/Q _09186_/B _11522_/S vssd1 vssd1 vccd1 vccd1 _11518_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12498_ _13243_/CLK _12498_/D vssd1 vssd1 vccd1 vccd1 _12498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11449_ _12924_/Q _10793_/A _11449_/S vssd1 vssd1 vccd1 vccd1 _11449_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13119_ _12168_/X _13119_/D _07181_/X vssd1 vssd1 vccd1 vccd1 _13119_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06990_ _06987_/Y _11882_/X _11879_/X _06989_/Y vssd1 vssd1 vccd1 vccd1 _06995_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_112_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08660_ _11927_/X _08654_/X _12718_/Q _08655_/X vssd1 vssd1 vccd1 vccd1 _12718_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07611_ _07611_/A vssd1 vssd1 vccd1 vccd1 _07611_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08591_ _08591_/A vssd1 vssd1 vccd1 vccd1 _08591_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07542_ _12996_/Q _07531_/X _09226_/A _07532_/X _07538_/X vssd1 vssd1 vccd1 vccd1
+ _12996_/D sky130_fd_sc_hd__o221a_1
XFILLER_201_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07473_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07473_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09212_ _12477_/Q _09207_/X _09242_/A _09208_/X vssd1 vssd1 vccd1 vccd1 _12477_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06424_ _10717_/A vssd1 vssd1 vccd1 vccd1 _06425_/A sky130_fd_sc_hd__inv_2
XFILLER_194_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09143_ _12504_/Q _09143_/B vssd1 vssd1 vccd1 vccd1 _09144_/B sky130_fd_sc_hd__or2_1
X_06355_ _08519_/A vssd1 vssd1 vccd1 vccd1 _08504_/A sky130_fd_sc_hd__buf_2
X_09074_ _09439_/A _10527_/D vssd1 vssd1 vccd1 vccd1 _09083_/A sky130_fd_sc_hd__or2_2
XFILLER_190_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06286_ _09009_/A vssd1 vssd1 vccd1 vccd1 _06416_/A sky130_fd_sc_hd__buf_6
XFILLER_147_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08025_ _08025_/A vssd1 vssd1 vccd1 vccd1 _08041_/A sky130_fd_sc_hd__inv_2
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09976_ _09981_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _10137_/A sky130_fd_sc_hd__or2_4
XFILLER_118_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08927_ _08927_/A _08927_/B vssd1 vssd1 vccd1 vccd1 _10636_/A sky130_fd_sc_hd__or2_1
XFILLER_29_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08858_ _08866_/A vssd1 vssd1 vccd1 vccd1 _08858_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07809_ _12924_/Q vssd1 vssd1 vccd1 vccd1 _07809_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08789_ _08789_/A vssd1 vssd1 vccd1 vccd1 _08789_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_73_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10820_ _10821_/B _10819_/X _10821_/B _10819_/X vssd1 vssd1 vccd1 vccd1 _12327_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_77_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_98_wb_clk_i _13219_/CLK vssd1 vssd1 vccd1 vccd1 _13193_/CLK sky130_fd_sc_hd__clkbuf_16
X_10751_ _11083_/A vssd1 vssd1 vccd1 vccd1 _10751_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12434_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10682_ _12445_/Q _12446_/Q _08946_/B vssd1 vssd1 vccd1 vccd1 _10682_/X sky130_fd_sc_hd__a21bo_1
XFILLER_41_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12421_ _12422_/CLK _12421_/D vssd1 vssd1 vccd1 vccd1 _12421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12352_ _12353_/CLK _12352_/D vssd1 vssd1 vccd1 vccd1 _12352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11303_ vssd1 vssd1 vccd1 vccd1 _11303_/HI _11303_/LO sky130_fd_sc_hd__conb_1
XFILLER_5_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12283_ _12296_/CLK _12283_/D vssd1 vssd1 vccd1 vccd1 _12283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11234_ vssd1 vssd1 vccd1 vccd1 _11234_/HI _11234_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11165_ vssd1 vssd1 vccd1 vccd1 _11165_/HI _11165_/LO sky130_fd_sc_hd__conb_1
XFILLER_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10116_ _12626_/Q vssd1 vssd1 vccd1 vccd1 _10116_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11096_ _10763_/X _11054_/A _06379_/X _11055_/A _11060_/X vssd1 vssd1 vccd1 vccd1
+ _11096_/X sky130_fd_sc_hd__a221o_1
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput340 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 input340/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput351 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 input351/X sky130_fd_sc_hd__clkbuf_2
Xinput362 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _09293_/B sky130_fd_sc_hd__buf_1
X_10047_ _10796_/A _10047_/B _10151_/A vssd1 vssd1 vccd1 vccd1 _11878_/S sky130_fd_sc_hd__and3_4
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11998_ _11061_/X _11056_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _11998_/X sky130_fd_sc_hd__mux2_2
XFILLER_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10949_ _12532_/Q _12344_/Q _12533_/Q _12345_/Q _10948_/X vssd1 vssd1 vccd1 vccd1
+ _10949_/X sky130_fd_sc_hd__a221o_1
XFILLER_17_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ _12619_/CLK _12619_/D vssd1 vssd1 vccd1 vccd1 _12619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06140_ _06067_/A _06067_/B _06067_/X _06064_/A vssd1 vssd1 vccd1 vccd1 _06140_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06071_ _12732_/Q _12700_/Q _12732_/Q _12700_/Q vssd1 vssd1 vccd1 vccd1 _06075_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_32_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09830_ _09770_/X _09868_/C _09825_/Y _09828_/X _09829_/X vssd1 vssd1 vccd1 vccd1
+ _09832_/B sky130_fd_sc_hd__o311a_1
XFILLER_112_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09761_ _09755_/Y _09760_/X _09755_/Y _09760_/X vssd1 vssd1 vccd1 vccd1 _09762_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_06973_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06973_/X sky130_fd_sc_hd__clkbuf_1
X_08712_ _08714_/A vssd1 vssd1 vccd1 vccd1 _08712_/X sky130_fd_sc_hd__clkbuf_1
X_09692_ _09687_/X _09691_/X _09687_/X _09691_/X vssd1 vssd1 vccd1 vccd1 _09692_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08643_ _08653_/A vssd1 vssd1 vccd1 vccd1 _08643_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_199_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _08715_/A vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__buf_2
XFILLER_82_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ _13002_/Q _07520_/Y _07568_/A _07520_/A _07522_/Y vssd1 vssd1 vccd1 vccd1
+ _13002_/D sky130_fd_sc_hd__o221a_1
XFILLER_23_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07456_ _07458_/A vssd1 vssd1 vccd1 vccd1 _07456_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06407_ _13240_/Q vssd1 vssd1 vccd1 vccd1 _06407_/X sky130_fd_sc_hd__buf_2
XFILLER_194_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07387_ _07391_/A vssd1 vssd1 vccd1 vccd1 _07387_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09126_ _12516_/Q _09123_/X _08005_/X _09124_/X vssd1 vssd1 vccd1 vccd1 _12516_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06338_ _06344_/A vssd1 vssd1 vccd1 vccd1 _06338_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09057_ _09058_/A _12149_/X vssd1 vssd1 vccd1 vccd1 _12560_/D sky130_fd_sc_hd__nor2b_1
X_06269_ _07742_/B vssd1 vssd1 vccd1 vccd1 _06269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08008_ _08018_/A vssd1 vssd1 vccd1 vccd1 _08008_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_117_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_145_wb_clk_i _12844_/CLK vssd1 vssd1 vccd1 vccd1 _12872_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09959_ _08753_/Y _09897_/A _06200_/X _09892_/A _09941_/A vssd1 vssd1 vccd1 vccd1
+ _09959_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12970_ _12984_/CLK _12970_/D vssd1 vssd1 vccd1 vccd1 _12970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11921_ _11920_/X _12442_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11921_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _11035_/X _10700_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _11852_/X sky130_fd_sc_hd__mux2_2
XPHY_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _12511_/Q _12323_/Q _10799_/Y _10801_/X vssd1 vssd1 vccd1 vccd1 _10806_/A
+ sky130_fd_sc_hd__a22o_1
XPHY_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _12120_/X _12480_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11783_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10734_ _10730_/X _10731_/X _06362_/X _10732_/X _10733_/X vssd1 vssd1 vccd1 vccd1
+ _10734_/X sky130_fd_sc_hd__a221o_1
XFILLER_201_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10665_ _08944_/A _08944_/B _09311_/A vssd1 vssd1 vccd1 vccd1 _10665_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ _12410_/CLK _12404_/D vssd1 vssd1 vccd1 vccd1 _12404_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10596_ _10603_/A _10595_/Y _09385_/Y _10526_/B vssd1 vssd1 vccd1 vccd1 _10607_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_154_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12335_ _12337_/CLK _12335_/D vssd1 vssd1 vccd1 vccd1 _12335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12266_ _12265_/X _12653_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12266_/X sky130_fd_sc_hd__mux2_2
XFILLER_141_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11217_ vssd1 vssd1 vccd1 vccd1 _11217_/HI _11217_/LO sky130_fd_sc_hd__conb_1
XFILLER_123_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12197_ _06583_/A _10744_/Y _12760_/Q vssd1 vssd1 vccd1 vccd1 _12198_/S sky130_fd_sc_hd__mux2_8
XFILLER_150_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11148_ vssd1 vssd1 vccd1 vccd1 _11148_/HI _11148_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11079_ _11079_/A vssd1 vssd1 vccd1 vccd1 _11079_/Y sky130_fd_sc_hd__inv_2
Xinput170 la_oenb[102] vssd1 vssd1 vccd1 vccd1 input170/X sky130_fd_sc_hd__buf_1
Xinput181 la_oenb[112] vssd1 vssd1 vccd1 vccd1 input181/X sky130_fd_sc_hd__buf_1
XFILLER_37_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput192 la_oenb[122] vssd1 vssd1 vccd1 vccd1 input192/X sky130_fd_sc_hd__buf_1
XFILLER_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07310_ _13075_/Q _07285_/A _07309_/X _07284_/A vssd1 vssd1 vccd1 vccd1 _13075_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08290_ _12831_/Q _11606_/X _08292_/S vssd1 vssd1 vccd1 vccd1 _12831_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07241_ _07251_/A vssd1 vssd1 vccd1 vccd1 _07241_/X sky130_fd_sc_hd__clkbuf_1
X_07172_ _11524_/X _07160_/X _13123_/Q _07161_/X vssd1 vssd1 vccd1 vccd1 _13123_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06123_ _06117_/Y _06118_/Y _06115_/Y _06116_/Y vssd1 vssd1 vccd1 vccd1 _06123_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_8_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput600 _12286_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_105_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06054_ _12705_/Q vssd1 vssd1 vccd1 vccd1 _06054_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09813_ _09810_/Y _09812_/Y _13226_/Q _09812_/A vssd1 vssd1 vccd1 vccd1 _09813_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09744_ _09742_/A _09742_/B _09743_/Y vssd1 vssd1 vccd1 vccd1 _09745_/B sky130_fd_sc_hd__a21o_1
X_06956_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06956_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09675_ _09675_/A _09714_/A vssd1 vssd1 vccd1 vccd1 _09675_/X sky130_fd_sc_hd__or2_1
X_06887_ _06887_/A vssd1 vssd1 vccd1 vccd1 _06887_/X sky130_fd_sc_hd__buf_2
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08626_ _11940_/X _08624_/X _12731_/Q _08625_/X vssd1 vssd1 vccd1 vccd1 _12731_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _12616_/D _08557_/B _08562_/B vssd1 vssd1 vccd1 vccd1 _08558_/S sky130_fd_sc_hd__or3_1
XFILLER_39_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07508_ _13006_/Q vssd1 vssd1 vccd1 vccd1 _07508_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08488_ _13064_/Q vssd1 vssd1 vccd1 vccd1 _08488_/Y sky130_fd_sc_hd__inv_2
XPHY_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07439_ _07443_/A vssd1 vssd1 vccd1 vccd1 _07439_/X sky130_fd_sc_hd__clkbuf_1
XPHY_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10450_ _10450_/A vssd1 vssd1 vccd1 vccd1 _10452_/B sky130_fd_sc_hd__inv_2
XFILLER_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09109_ _12529_/Q _09107_/X input339/X _09108_/X vssd1 vssd1 vccd1 vccd1 _12529_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10381_ _10381_/A vssd1 vssd1 vccd1 vccd1 _10385_/C sky130_fd_sc_hd__inv_2
XFILLER_164_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12120_ _12119_/X _12436_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12120_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12051_ _11130_/X _11127_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _12051_/X sky130_fd_sc_hd__mux2_2
XFILLER_78_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11002_ _10988_/Y _10995_/Y _10990_/X _11001_/X vssd1 vssd1 vccd1 vccd1 _11002_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_133_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12953_ _12957_/CLK _12953_/D vssd1 vssd1 vccd1 vccd1 _12953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11904_ _08928_/A _10640_/Y _12321_/Q vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12974_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12884_ _12886_/CLK _12884_/D _08002_/X vssd1 vssd1 vccd1 vccd1 _12884_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _09942_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11835_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11766_ _11765_/X _12107_/X _11774_/S vssd1 vssd1 vccd1 vccd1 _12431_/D sky130_fd_sc_hd__mux2_1
XPHY_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10717_ _10717_/A vssd1 vssd1 vccd1 vccd1 _10717_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11697_ _11399_/X _09180_/D _11703_/S vssd1 vssd1 vccd1 vccd1 _11697_/X sky130_fd_sc_hd__mux2_1
XPHY_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10648_ _11906_/X vssd1 vssd1 vccd1 vccd1 _10648_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10579_ _10579_/A _10579_/B vssd1 vssd1 vccd1 vccd1 _10579_/X sky130_fd_sc_hd__or2_1
XFILLER_6_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12318_ _12987_/CLK _12318_/D vssd1 vssd1 vccd1 vccd1 _12318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12249_ _12779_/Q _12852_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12249_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06810_ _06860_/A _06861_/B vssd1 vssd1 vccd1 vccd1 _06810_/Y sky130_fd_sc_hd__nand2_1
X_07790_ _09019_/B _07519_/B _11982_/S _12925_/Q vssd1 vssd1 vccd1 vccd1 _07790_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_7_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06741_ _06734_/A _06734_/B _06734_/X vssd1 vssd1 vccd1 vccd1 _06741_/X sky130_fd_sc_hd__a21bo_1
X_09460_ _12971_/Q _09440_/A _12605_/Q _07519_/B vssd1 vssd1 vccd1 vccd1 _09460_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06672_ _12046_/X vssd1 vssd1 vccd1 vccd1 _06672_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08411_ _12784_/Q _08401_/X _07986_/X _08403_/X vssd1 vssd1 vccd1 vccd1 _12784_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09391_ _12547_/Q _10610_/B _12452_/Q _09390_/Y vssd1 vssd1 vccd1 vccd1 _09391_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08342_ _08352_/A vssd1 vssd1 vccd1 vccd1 _08342_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08273_ _13076_/Q vssd1 vssd1 vccd1 vccd1 _08273_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07224_ _07236_/A vssd1 vssd1 vccd1 vccd1 _07224_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07155_ _07167_/A vssd1 vssd1 vccd1 vccd1 _07155_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_145_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06106_ _12691_/Q vssd1 vssd1 vccd1 vccd1 _06106_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07086_ _09267_/C vssd1 vssd1 vccd1 vccd1 _09073_/A sky130_fd_sc_hd__inv_2
XFILLER_191_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput430 _11210_/LO vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__clkbuf_2
Xoutput441 _11186_/LO vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_69_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput452 _11321_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06037_ _06037_/A vssd1 vssd1 vccd1 vccd1 _06046_/A sky130_fd_sc_hd__inv_2
Xoutput463 _11331_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__clkbuf_2
Xoutput474 _11341_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__clkbuf_2
Xoutput485 _11217_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput496 _11218_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07988_ _08038_/A vssd1 vssd1 vccd1 vccd1 _08004_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09727_ _09722_/X _09726_/X _09722_/X _09726_/X vssd1 vssd1 vccd1 vccd1 _09727_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_132_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06939_ _13182_/Q vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__inv_2
XFILLER_132_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09658_ _09641_/A _09657_/A _09641_/Y _09657_/Y vssd1 vssd1 vccd1 vccd1 _09673_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08609_ _08716_/A vssd1 vssd1 vccd1 vccd1 _08686_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_163_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09589_/A vssd1 vssd1 vccd1 vccd1 _09589_/Y sky130_fd_sc_hd__inv_2
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _10490_/X _12987_/Q _12307_/D vssd1 vssd1 vccd1 vccd1 _11620_/X sky130_fd_sc_hd__mux2_1
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _12808_/Q _09186_/A _11558_/S vssd1 vssd1 vccd1 vccd1 _11551_/X sky130_fd_sc_hd__mux2_1
XPHY_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10502_ _12507_/Q _09146_/B _09147_/B vssd1 vssd1 vccd1 vccd1 _10502_/X sky130_fd_sc_hd__a21bo_1
XPHY_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11482_ _10317_/Y _09184_/A _11487_/S vssd1 vssd1 vccd1 vccd1 _11482_/X sky130_fd_sc_hd__mux2_1
XPHY_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_160_wb_clk_i clkbuf_opt_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _12540_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13221_ _13223_/CLK _13221_/D _06575_/X vssd1 vssd1 vccd1 vccd1 _13221_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10433_ _10433_/A _10433_/B _10433_/C vssd1 vssd1 vccd1 vccd1 _10439_/C sky130_fd_sc_hd__or3_4
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13152_ _13152_/CLK _13152_/D _07068_/X vssd1 vssd1 vccd1 vccd1 _13152_/Q sky130_fd_sc_hd__dfrtp_4
X_10364_ _10362_/B _10368_/D _10368_/A vssd1 vssd1 vccd1 vccd1 _10365_/C sky130_fd_sc_hd__o21a_1
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ _12102_/X _12430_/Q _12103_/S vssd1 vssd1 vccd1 vccd1 _12103_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13083_ _12167_/X _13083_/D _07278_/X vssd1 vssd1 vccd1 vccd1 _13083_/Q sky130_fd_sc_hd__dfrtp_1
X_10295_ _13269_/Q vssd1 vssd1 vccd1 vccd1 _10295_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12034_ _11094_/X _11089_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _12034_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12936_ _12937_/CLK _12936_/D vssd1 vssd1 vccd1 vccd1 _12936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12867_ _12870_/CLK _12867_/D _08047_/X vssd1 vssd1 vccd1 vccd1 _12867_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11818_ _12096_/X _11817_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11818_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12798_ _12892_/CLK _12798_/D _08370_/X vssd1 vssd1 vccd1 vccd1 _12798_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11749_ _11374_/X _11748_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11749_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08960_ _08962_/A vssd1 vssd1 vccd1 vccd1 _08960_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07911_ _07917_/A vssd1 vssd1 vccd1 vccd1 _07911_/X sky130_fd_sc_hd__clkbuf_1
X_08891_ _08883_/X _06300_/Y _08878_/X _12632_/Q vssd1 vssd1 vccd1 vccd1 _12632_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_29_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07842_ _07842_/A _07842_/B _07836_/X _07841_/X vssd1 vssd1 vccd1 vccd1 _07880_/B
+ sky130_fd_sc_hd__or4bb_4
XFILLER_116_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07773_ _12935_/Q _11648_/S _12936_/Q _07769_/X _07569_/X vssd1 vssd1 vccd1 vccd1
+ _12936_/D sky130_fd_sc_hd__a221o_1
XFILLER_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09512_ _13171_/Q vssd1 vssd1 vccd1 vccd1 _09526_/B sky130_fd_sc_hd__inv_2
X_06724_ _12033_/X _06724_/B vssd1 vssd1 vccd1 vccd1 _06724_/X sky130_fd_sc_hd__or2_1
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09443_ _09443_/A vssd1 vssd1 vccd1 vccd1 _09451_/A sky130_fd_sc_hd__inv_2
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06655_ _06507_/X _06651_/Y _06608_/X _06654_/X vssd1 vssd1 vccd1 vccd1 _13214_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09374_ _12542_/Q vssd1 vssd1 vccd1 vccd1 _09374_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06586_ _06586_/A vssd1 vssd1 vccd1 vccd1 _06587_/B sky130_fd_sc_hd__inv_2
XFILLER_33_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08325_ _08325_/A vssd1 vssd1 vccd1 vccd1 _08325_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_178_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08256_ _07293_/X _08251_/X _07406_/X vssd1 vssd1 vccd1 vccd1 _12841_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07207_ _11577_/X _07201_/X _13112_/Q _07204_/X vssd1 vssd1 vccd1 vccd1 _13112_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08187_ _10439_/B vssd1 vssd1 vccd1 vccd1 _08187_/X sky130_fd_sc_hd__buf_1
XFILLER_119_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07138_ _11537_/X _07130_/X _13136_/Q _07131_/X vssd1 vssd1 vccd1 vccd1 _13136_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07069_ _07069_/A vssd1 vssd1 vccd1 vccd1 _07069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10080_ _10078_/Y _10023_/X _10079_/Y _10025_/X vssd1 vssd1 vccd1 vccd1 _10088_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_88_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10982_ _12539_/Q _12351_/Q _12539_/Q _12351_/Q vssd1 vssd1 vccd1 vccd1 _11000_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12721_ _13162_/CLK _12721_/D _08649_/X vssd1 vssd1 vccd1 vccd1 _12721_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _13159_/CLK _12652_/D _08840_/X vssd1 vssd1 vccd1 vccd1 _12652_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_169_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _10471_/X _10792_/B _11603_/S vssd1 vssd1 vccd1 vccd1 _11603_/X sky130_fd_sc_hd__mux2_1
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ _12586_/CLK _12583_/D vssd1 vssd1 vccd1 vccd1 _12583_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11534_ _12823_/Q _09180_/C _11543_/S vssd1 vssd1 vccd1 vccd1 _11534_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11465_ _12908_/Q _10528_/B _11469_/S vssd1 vssd1 vccd1 vccd1 _11465_/X sky130_fd_sc_hd__mux2_1
X_13204_ _13205_/CLK _13204_/D _06738_/X vssd1 vssd1 vccd1 vccd1 _13204_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10416_ _10418_/B vssd1 vssd1 vccd1 vccd1 _10416_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11396_ _10622_/X _12414_/D _11889_/S vssd1 vssd1 vccd1 vccd1 _11396_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13135_ _12168_/X _13135_/D _07140_/X vssd1 vssd1 vccd1 vccd1 _13135_/Q sky130_fd_sc_hd__dfrtp_1
X_10347_ _10352_/C vssd1 vssd1 vccd1 vccd1 _10349_/B sky130_fd_sc_hd__inv_2
XFILLER_174_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13066_ _12165_/X _13066_/D _07341_/X vssd1 vssd1 vccd1 vccd1 _13066_/Q sky130_fd_sc_hd__dfrtp_1
X_10278_ _13094_/Q _10276_/X _13126_/Q _10277_/X vssd1 vssd1 vccd1 vccd1 _10278_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12017_ _11066_/X _11059_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12017_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12919_ _12166_/X _12919_/D _07903_/X vssd1 vssd1 vccd1 vccd1 _12919_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06440_ _06658_/A vssd1 vssd1 vccd1 vccd1 _06440_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06371_ _13250_/Q vssd1 vssd1 vccd1 vccd1 _06371_/X sky130_fd_sc_hd__buf_2
XFILLER_187_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08110_ _08107_/Y _10484_/A _08109_/Y _12806_/Q vssd1 vssd1 vccd1 vccd1 _08110_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09090_ _09123_/A vssd1 vssd1 vccd1 vccd1 _09124_/A sky130_fd_sc_hd__inv_2
XFILLER_30_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08041_ _08041_/A vssd1 vssd1 vccd1 vccd1 _08041_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09992_ _08794_/Y _09968_/X _06263_/Y _09972_/X _09991_/X vssd1 vssd1 vccd1 vccd1
+ _09992_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_89_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08943_ _12427_/Q _11370_/S vssd1 vssd1 vccd1 vccd1 _08944_/B sky130_fd_sc_hd__and2b_1
XFILLER_9_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08874_ _07747_/X _06351_/X _08837_/A _12638_/Q vssd1 vssd1 vccd1 vccd1 _12638_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07825_ _13011_/Q _07823_/Y _13034_/Q _07824_/Y vssd1 vssd1 vccd1 vccd1 _07825_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07756_ _12582_/Q _07756_/B vssd1 vssd1 vccd1 vccd1 _07757_/B sky130_fd_sc_hd__or2_1
X_06707_ _06707_/A vssd1 vssd1 vccd1 vccd1 _13208_/D sky130_fd_sc_hd__inv_2
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07687_ _12964_/Q _07682_/A _07682_/Y _07686_/X _09283_/A vssd1 vssd1 vccd1 vccd1
+ _12964_/D sky130_fd_sc_hd__a221o_1
XFILLER_73_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09426_ _12461_/Q _09423_/Y _12465_/Q _10579_/A _09425_/X vssd1 vssd1 vccd1 vccd1
+ _09426_/X sky130_fd_sc_hd__o221a_1
XFILLER_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06638_ _06356_/X _07019_/A _06427_/X _11071_/A _06637_/Y vssd1 vssd1 vccd1 vccd1
+ _10765_/A sky130_fd_sc_hd__o221a_2
XFILLER_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09357_ _12547_/Q vssd1 vssd1 vccd1 vccd1 _09357_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06569_ _06569_/A vssd1 vssd1 vccd1 vccd1 _06573_/A sky130_fd_sc_hd__inv_2
XFILLER_200_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08308_ _08311_/A vssd1 vssd1 vccd1 vccd1 _08308_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_100_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09288_ _09288_/A _09288_/B vssd1 vssd1 vccd1 vccd1 _09288_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08239_ _13087_/Q vssd1 vssd1 vccd1 vccd1 _08239_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11250_ vssd1 vssd1 vccd1 vccd1 _11250_/HI _11250_/LO sky130_fd_sc_hd__conb_1
XFILLER_134_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10201_ _12630_/Q vssd1 vssd1 vccd1 vccd1 _10201_/Y sky130_fd_sc_hd__inv_2
X_11181_ vssd1 vssd1 vccd1 vccd1 _11181_/HI _11181_/LO sky130_fd_sc_hd__conb_1
XFILLER_69_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10132_ _13013_/Q _10276_/A _13046_/Q _10277_/A vssd1 vssd1 vccd1 vccd1 _10132_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10063_ _13256_/Q vssd1 vssd1 vccd1 vccd1 _10063_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10965_ _12534_/Q _12346_/Q _10958_/Y vssd1 vssd1 vccd1 vccd1 _10965_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ _12707_/CLK _12704_/D _08693_/X vssd1 vssd1 vccd1 vccd1 _12704_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10896_ _10921_/A vssd1 vssd1 vccd1 vccd1 _10896_/Y sky130_fd_sc_hd__inv_2
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12635_ _13158_/CLK _12635_/D _08882_/X vssd1 vssd1 vccd1 vccd1 _12635_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12566_ _12570_/CLK _12566_/D vssd1 vssd1 vccd1 vccd1 _12566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ _12806_/Q _09185_/C _11546_/S vssd1 vssd1 vccd1 vccd1 _11517_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12497_ _13243_/CLK _12497_/D vssd1 vssd1 vccd1 vccd1 _12497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11448_ _12923_/Q _10793_/B _11449_/S vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11379_ _10570_/Y _12398_/D _11392_/S vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13118_ _12168_/X _13118_/D _07183_/X vssd1 vssd1 vccd1 vccd1 _13118_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_79_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13049_ _12165_/X _13049_/D _07383_/X vssd1 vssd1 vccd1 vccd1 _13049_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07610_ _07610_/A vssd1 vssd1 vccd1 vccd1 _07610_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08590_ _11953_/X _08575_/X _12744_/Q _08578_/X vssd1 vssd1 vccd1 vccd1 _12744_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07541_ _12997_/Q _07531_/X _07562_/A _07532_/X _07538_/X vssd1 vssd1 vccd1 vccd1
+ _12997_/D sky130_fd_sc_hd__o221a_1
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07472_ _11458_/X _07459_/X _13017_/Q _07460_/X vssd1 vssd1 vccd1 vccd1 _13017_/D
+ sky130_fd_sc_hd__a22o_1
X_09211_ _12478_/Q _09207_/X _09243_/D _09208_/X vssd1 vssd1 vccd1 vccd1 _12478_/D
+ sky130_fd_sc_hd__a22o_1
X_06423_ _10714_/A _10714_/B _12770_/Q vssd1 vssd1 vccd1 vccd1 _10717_/A sky130_fd_sc_hd__o21ai_4
XFILLER_72_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09142_ _12503_/Q _09142_/B vssd1 vssd1 vccd1 vccd1 _09143_/B sky130_fd_sc_hd__or2_1
XFILLER_33_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06354_ _12945_/Q vssd1 vssd1 vccd1 vccd1 _08519_/A sky130_fd_sc_hd__inv_2
XFILLER_175_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09073_ _09073_/A _11030_/B vssd1 vssd1 vccd1 vccd1 _10527_/D sky130_fd_sc_hd__or2_4
X_06285_ _08854_/A vssd1 vssd1 vccd1 vccd1 _09009_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08024_ _08040_/A vssd1 vssd1 vccd1 vccd1 _08024_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09975_ _12860_/Q vssd1 vssd1 vccd1 vccd1 _09975_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08926_ _08926_/A _08926_/B vssd1 vssd1 vccd1 vccd1 _08927_/B sky130_fd_sc_hd__or2_1
XFILLER_103_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08857_ _08849_/X _06311_/Y _08852_/X _12646_/Q vssd1 vssd1 vccd1 vccd1 _12646_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07808_ _13019_/Q vssd1 vssd1 vccd1 vccd1 _07808_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08788_ _08787_/Y _08781_/X _06255_/X _08764_/A vssd1 vssd1 vccd1 vccd1 _12672_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07739_ _07749_/A vssd1 vssd1 vccd1 vccd1 _07739_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10750_ _11075_/A vssd1 vssd1 vccd1 vccd1 _10750_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09409_ _12459_/Q _09394_/A _12547_/Q _10610_/B vssd1 vssd1 vccd1 vccd1 _09409_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10681_ _12445_/Q _12090_/S _10680_/Y _09318_/A vssd1 vssd1 vccd1 vccd1 _10681_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_179_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12420_ _12422_/CLK _12420_/D vssd1 vssd1 vccd1 vccd1 _12420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12351_ _12353_/CLK _12351_/D vssd1 vssd1 vccd1 vccd1 _12351_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_67_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12975_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ vssd1 vssd1 vccd1 vccd1 _11302_/HI _11302_/LO sky130_fd_sc_hd__conb_1
XFILLER_153_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _10314_/X _12908_/Q _11878_/X _10312_/Y _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12298_/D sky130_fd_sc_hd__mux4_2
XFILLER_154_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11233_ vssd1 vssd1 vccd1 vccd1 _11233_/HI _11233_/LO sky130_fd_sc_hd__conb_1
XFILLER_122_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11164_ vssd1 vssd1 vccd1 vccd1 _11164_/HI _11164_/LO sky130_fd_sc_hd__conb_1
XFILLER_136_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10115_ _07799_/Y _10070_/X _10114_/X vssd1 vssd1 vccd1 vccd1 _10115_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11095_ _10755_/X _11071_/X _13250_/Q _11058_/X _11072_/X vssd1 vssd1 vccd1 vccd1
+ _11095_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput330 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 _07993_/A sky130_fd_sc_hd__buf_2
XFILLER_96_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput341 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 input341/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput352 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 _10793_/B sky130_fd_sc_hd__buf_4
X_10046_ _10113_/A vssd1 vssd1 vccd1 vccd1 _10047_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_76_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput363 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _09293_/C sky130_fd_sc_hd__buf_1
XFILLER_17_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11997_ _11076_/X _11068_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _11997_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10948_ _10930_/Y _10946_/X _10947_/Y _12532_/Q _12344_/Q vssd1 vssd1 vccd1 vccd1
+ _10948_/X sky130_fd_sc_hd__o32a_1
XFILLER_32_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10879_ _12524_/Q vssd1 vssd1 vccd1 vccd1 _10879_/Y sky130_fd_sc_hd__inv_2
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12618_ _13241_/CLK _12618_/D _08959_/X vssd1 vssd1 vccd1 vccd1 _12618_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12549_ _12875_/CLK _12549_/D _09069_/X vssd1 vssd1 vccd1 vccd1 _12549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_129_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06070_ _06172_/B _06182_/B vssd1 vssd1 vccd1 vccd1 _06070_/X sky130_fd_sc_hd__or2_1
XFILLER_172_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09760_ _09756_/X _09759_/X _09756_/X _09759_/X vssd1 vssd1 vccd1 vccd1 _09760_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06972_ _06457_/X _09578_/B _06459_/X _06971_/Y vssd1 vssd1 vccd1 vccd1 _13179_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_140_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08711_ _11831_/X _08700_/X _12697_/Q _08701_/X vssd1 vssd1 vccd1 vccd1 _12697_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09691_ _13203_/Q _09690_/A _09689_/Y _09690_/Y vssd1 vssd1 vccd1 vccd1 _09691_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_6_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08642_ _08642_/A vssd1 vssd1 vccd1 vccd1 _08653_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _12616_/Q _09469_/A vssd1 vssd1 vccd1 vccd1 _08715_/A sky130_fd_sc_hd__or2_2
XPHY_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07524_ _13003_/Q _07520_/Y _09226_/B _07520_/A _07522_/Y vssd1 vssd1 vccd1 vccd1
+ _13003_/D sky130_fd_sc_hd__o221a_1
XPHY_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07455_ _11465_/X _07444_/X _13024_/Q _07445_/X vssd1 vssd1 vccd1 vccd1 _13024_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06406_ _06412_/A vssd1 vssd1 vccd1 vccd1 _06406_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07386_ _11425_/X _07384_/X _13049_/Q _07385_/X vssd1 vssd1 vccd1 vccd1 _13049_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09125_ _12517_/Q _09123_/X _07545_/X _09124_/X vssd1 vssd1 vccd1 vccd1 _12517_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06337_ _07742_/B _06314_/X _06336_/Y _13258_/Q _06306_/A vssd1 vssd1 vccd1 vccd1
+ _13258_/D sky130_fd_sc_hd__a32o_1
XFILLER_163_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ _09058_/A _12150_/X vssd1 vssd1 vccd1 vccd1 _12561_/D sky130_fd_sc_hd__nor2b_1
X_06268_ _12608_/Q vssd1 vssd1 vccd1 vccd1 _07742_/B sky130_fd_sc_hd__clkbuf_2
X_08007_ _08038_/A vssd1 vssd1 vccd1 vccd1 _08018_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06199_ _06026_/Y _06027_/Y _06030_/A _06198_/X vssd1 vssd1 vccd1 vccd1 _06199_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_1_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09958_ _08756_/Y _09952_/X _06204_/X _09892_/A _09941_/A vssd1 vssd1 vccd1 vccd1
+ _09958_/Y sky130_fd_sc_hd__o221ai_2
X_08909_ _08898_/X _06336_/Y _08908_/X _12625_/Q vssd1 vssd1 vccd1 vccd1 _12625_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_170_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09889_ _12654_/Q _12611_/Q _06351_/X _09547_/A _09888_/Y vssd1 vssd1 vccd1 vccd1
+ _09889_/X sky130_fd_sc_hd__a221o_1
XFILLER_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11920_ _12442_/Q _11919_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _11920_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _09962_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11851_/X sky130_fd_sc_hd__mux2_1
XPHY_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _10799_/Y _10801_/X _10799_/Y _10801_/X vssd1 vssd1 vccd1 vccd1 _12323_/D
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _11781_/X _12136_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12435_/D sky130_fd_sc_hd__mux2_1
XPHY_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ _12116_/X vssd1 vssd1 vccd1 vccd1 _10733_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10664_ _08944_/B _10663_/X _09311_/A vssd1 vssd1 vccd1 vccd1 _10664_/X sky130_fd_sc_hd__o21a_1
XFILLER_186_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12403_ _12410_/CLK _12403_/D vssd1 vssd1 vccd1 vccd1 _12403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10595_ _12407_/D _10594_/A _12408_/D vssd1 vssd1 vccd1 vccd1 _10595_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_154_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12334_ _12802_/CLK _12334_/D vssd1 vssd1 vccd1 vccd1 _12334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12265_ _12787_/Q _12860_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12265_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11216_ vssd1 vssd1 vccd1 vccd1 _11216_/HI _11216_/LO sky130_fd_sc_hd__conb_1
X_12196_ _10753_/X _10756_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _12196_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11147_ _11147_/A vssd1 vssd1 vccd1 vccd1 _11147_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11078_ _10696_/X _11077_/X _06404_/X _10760_/X _10761_/X vssd1 vssd1 vccd1 vccd1
+ _11078_/X sky130_fd_sc_hd__a221o_1
Xinput160 la_data_in[94] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_hd__buf_1
Xinput171 la_oenb[103] vssd1 vssd1 vccd1 vccd1 input171/X sky130_fd_sc_hd__buf_1
Xinput182 la_oenb[113] vssd1 vssd1 vccd1 vccd1 input182/X sky130_fd_sc_hd__buf_1
X_10029_ _12654_/Q vssd1 vssd1 vccd1 vccd1 _10029_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput193 la_oenb[123] vssd1 vssd1 vccd1 vccd1 input193/X sky130_fd_sc_hd__buf_1
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07240_ _11564_/X _07233_/X _13099_/Q _07234_/X vssd1 vssd1 vccd1 vccd1 _13099_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07171_ _07183_/A vssd1 vssd1 vccd1 vccd1 _07171_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06122_ _06122_/A _06122_/B vssd1 vssd1 vccd1 vccd1 _06122_/Y sky130_fd_sc_hd__nand2_2
Xoutput601 _12287_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__clkbuf_2
X_06053_ _12737_/Q vssd1 vssd1 vccd1 vccd1 _06053_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09812_ _09812_/A vssd1 vssd1 vccd1 vccd1 _09812_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09743_ _09743_/A vssd1 vssd1 vccd1 vccd1 _09743_/Y sky130_fd_sc_hd__inv_2
X_06955_ _06528_/X _06949_/X _06954_/Y _06841_/X _13180_/Q vssd1 vssd1 vccd1 vccd1
+ _13180_/D sky130_fd_sc_hd__a32o_1
XFILLER_100_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09674_ _09641_/Y _09659_/A _09657_/Y vssd1 vssd1 vccd1 vccd1 _09674_/Y sky130_fd_sc_hd__o21ai_1
X_06886_ _06886_/A vssd1 vssd1 vccd1 vccd1 _06886_/X sky130_fd_sc_hd__buf_2
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08625_ _08686_/A vssd1 vssd1 vccd1 vccd1 _08625_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _12609_/Q _08556_/B _08740_/A _08556_/D vssd1 vssd1 vccd1 vccd1 _08557_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_74_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07507_ _09185_/B vssd1 vssd1 vccd1 vccd1 _09228_/B sky130_fd_sc_hd__inv_2
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08487_ _13048_/Q _10333_/A _08485_/Y _12907_/Q _08486_/X vssd1 vssd1 vccd1 vccd1
+ _08493_/B sky130_fd_sc_hd__o221a_1
XPHY_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07438_ _11472_/X _07429_/X _13031_/Q _07430_/X vssd1 vssd1 vccd1 vccd1 _13031_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07369_ _07369_/A vssd1 vssd1 vccd1 vccd1 _07369_/X sky130_fd_sc_hd__buf_2
XFILLER_109_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09108_ _09116_/A vssd1 vssd1 vccd1 vccd1 _09108_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10380_ _10380_/A _10380_/B _10380_/C vssd1 vssd1 vccd1 vccd1 _10381_/A sky130_fd_sc_hd__or3_4
XFILLER_164_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09039_ _12571_/Q _09037_/X _08996_/D _09038_/Y vssd1 vssd1 vccd1 vccd1 _12571_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12050_ _10749_/X _11123_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _12050_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11001_ _12540_/Q _12352_/Q _10993_/X _12541_/Q _12353_/Q vssd1 vssd1 vccd1 vccd1
+ _11001_/X sky130_fd_sc_hd__a32o_1
XFILLER_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12952_ _12957_/CLK _12952_/D vssd1 vssd1 vccd1 vccd1 _12952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11903_ _08927_/A _10637_/X _12321_/Q vssd1 vssd1 vccd1 vccd1 _11903_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12883_ _12886_/CLK _12883_/D _08004_/X vssd1 vssd1 vccd1 vccd1 _12883_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _09936_/Y _12859_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11834_/X sky130_fd_sc_hd__mux2_1
XPHY_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _12107_/X _11764_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_82_wb_clk_i _12960_/CLK vssd1 vssd1 vccd1 vccd1 _13252_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_201_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _13243_/Q vssd1 vssd1 vccd1 vccd1 _11033_/A sky130_fd_sc_hd__inv_2
XFILLER_9_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _11695_/X _11402_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12390_/D sky130_fd_sc_hd__mux2_1
XPHY_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10647_ _12423_/Q _10643_/Y _08931_/A vssd1 vssd1 vccd1 vccd1 _10647_/Y sky130_fd_sc_hd__o21ai_1
X_10578_ _10579_/B vssd1 vssd1 vccd1 vccd1 _10578_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12317_ _12999_/CLK _12317_/D vssd1 vssd1 vccd1 vccd1 _12317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12248_ _12247_/X _12644_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12248_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12179_ _11144_/X _11140_/X _12193_/S vssd1 vssd1 vccd1 vccd1 _12179_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06740_ _06725_/X _06729_/X _06730_/X vssd1 vssd1 vccd1 vccd1 _06740_/X sky130_fd_sc_hd__a21bo_1
XFILLER_77_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06671_ _06671_/A vssd1 vssd1 vccd1 vccd1 _06671_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08410_ _08420_/A vssd1 vssd1 vccd1 vccd1 _08410_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_184_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09390_ _12404_/D vssd1 vssd1 vccd1 vccd1 _09390_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08341_ _08372_/A vssd1 vssd1 vccd1 vccd1 _08352_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_177_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08272_ _13075_/Q vssd1 vssd1 vccd1 vccd1 _08272_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07223_ _07253_/A vssd1 vssd1 vccd1 vccd1 _07236_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07154_ _07154_/A vssd1 vssd1 vccd1 vccd1 _07167_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06105_ _12723_/Q vssd1 vssd1 vccd1 vccd1 _06105_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07085_ _07547_/A vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__buf_2
Xoutput420 _11201_/LO vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput431 _11211_/LO vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__clkbuf_2
XFILLER_191_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput442 _11187_/LO vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__clkbuf_2
X_06036_ _12744_/Q _12712_/Q _12744_/Q _12712_/Q vssd1 vssd1 vccd1 vccd1 _06037_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput453 _11322_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__clkbuf_2
XFILLER_121_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput464 _11332_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__clkbuf_2
Xoutput475 _11342_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__clkbuf_2
Xoutput486 _11236_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__clkbuf_2
Xoutput497 _11246_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07987_ _12889_/Q _07974_/X _07986_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _12889_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09726_ _13209_/Q _09725_/A _09724_/Y _09725_/Y vssd1 vssd1 vccd1 vccd1 _09726_/X
+ sky130_fd_sc_hd__a22o_1
X_06938_ _06938_/A _06938_/B vssd1 vssd1 vccd1 vccd1 _06938_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09657_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09657_/Y sky130_fd_sc_hd__inv_2
X_06869_ _06916_/A vssd1 vssd1 vccd1 vccd1 _06869_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08608_ _08685_/A vssd1 vssd1 vccd1 vccd1 _08608_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09588_ _13184_/Q _13183_/Q _09604_/A _09604_/B vssd1 vssd1 vccd1 vccd1 _09589_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08539_ _08569_/A vssd1 vssd1 vccd1 vccd1 _08539_/X sky130_fd_sc_hd__clkbuf_1
XPHY_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _12807_/Q _09186_/B _11550_/S vssd1 vssd1 vccd1 vccd1 _11550_/X sky130_fd_sc_hd__mux2_1
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ _12506_/Q _09145_/B _09146_/B vssd1 vssd1 vccd1 vccd1 _10501_/X sky130_fd_sc_hd__a21bo_1
XPHY_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11481_ _12924_/Q _10793_/A _11481_/S vssd1 vssd1 vccd1 vccd1 _11481_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ _13227_/CLK _13220_/D _06580_/X vssd1 vssd1 vccd1 vccd1 _13220_/Q sky130_fd_sc_hd__dfrtp_1
X_10432_ _12814_/Q _10431_/B _10433_/B _10433_/C _10407_/X vssd1 vssd1 vccd1 vccd1
+ _10432_/X sky130_fd_sc_hd__o221a_1
XFILLER_183_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13151_ _13152_/CLK _13151_/D _07071_/X vssd1 vssd1 vccd1 vccd1 _13151_/Q sky130_fd_sc_hd__dfrtp_1
X_10363_ _10363_/A vssd1 vssd1 vccd1 vccd1 _10365_/B sky130_fd_sc_hd__inv_2
XFILLER_100_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12102_ _12430_/Q _12101_/X _12141_/S vssd1 vssd1 vccd1 vccd1 _12102_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13082_ _12167_/X _13082_/D _07280_/X vssd1 vssd1 vccd1 vccd1 _13082_/Q sky130_fd_sc_hd__dfrtp_4
X_10294_ _13022_/Q _10276_/X _13055_/Q _10277_/X vssd1 vssd1 vccd1 vccd1 _10294_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12033_ _11115_/X _11103_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12033_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12935_ _12973_/CLK _12935_/D vssd1 vssd1 vccd1 vccd1 _12935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _12868_/CLK _12866_/D _08049_/X vssd1 vssd1 vccd1 vccd1 _12866_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11817_ _09179_/C _11816_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11817_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12864_/CLK _12797_/D _08373_/X vssd1 vssd1 vccd1 vccd1 _12797_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_187_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11748_ _09185_/C _11747_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11748_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11679_ _11380_/X _09243_/D _11691_/S vssd1 vssd1 vccd1 vccd1 _11679_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07910_ _12917_/Q _11506_/X _07918_/S vssd1 vssd1 vccd1 vccd1 _12917_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08890_ _08897_/A vssd1 vssd1 vccd1 vccd1 _08890_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07841_ _13009_/Q _07822_/Y _13029_/Q _10373_/A _07840_/X vssd1 vssd1 vccd1 vccd1
+ _07841_/X sky130_fd_sc_hd__o221a_1
XFILLER_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07772_ _12578_/Q _11648_/S _12937_/Q _07769_/X _07569_/X vssd1 vssd1 vccd1 vccd1
+ _12937_/D sky130_fd_sc_hd__a221o_1
X_06723_ _12032_/X vssd1 vssd1 vccd1 vccd1 _06724_/B sky130_fd_sc_hd__inv_2
XFILLER_17_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09511_ _13172_/Q vssd1 vssd1 vccd1 vccd1 _09526_/A sky130_fd_sc_hd__inv_2
X_09442_ _09442_/A vssd1 vssd1 vccd1 vccd1 _09442_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06654_ _06645_/X _06632_/X _06652_/X _06653_/X vssd1 vssd1 vccd1 vccd1 _06654_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09373_ _09354_/Y _12400_/Q _09357_/Y _12416_/Q vssd1 vssd1 vccd1 vccd1 _09382_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06585_ _06427_/A _10745_/A _13254_/Q _07007_/A _11899_/X vssd1 vssd1 vccd1 vccd1
+ _06586_/A sky130_fd_sc_hd__a221o_2
XFILLER_75_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08324_ _12817_/Q _11592_/X _08335_/S vssd1 vssd1 vccd1 vccd1 _12817_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08255_ _08257_/A vssd1 vssd1 vccd1 vccd1 _08255_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07206_ _07206_/A vssd1 vssd1 vccd1 vccd1 _07206_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_192_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08186_ _12816_/Q vssd1 vssd1 vccd1 vccd1 _10439_/B sky130_fd_sc_hd__inv_2
XFILLER_119_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07137_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07137_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07068_ _07078_/A vssd1 vssd1 vccd1 vccd1 _07068_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_161_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06019_ _11726_/X _08562_/B vssd1 vssd1 vccd1 vccd1 _06272_/A sky130_fd_sc_hd__or2_2
XFILLER_87_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09709_ _09709_/A vssd1 vssd1 vccd1 vccd1 _09709_/Y sky130_fd_sc_hd__inv_2
X_10981_ _10975_/Y _10980_/Y _10975_/Y _10980_/Y vssd1 vssd1 vccd1 vccd1 _12350_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12720_ _13162_/CLK _12720_/D _08651_/X vssd1 vssd1 vccd1 vccd1 _12720_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_71_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ _12653_/CLK _12651_/D _08842_/X vssd1 vssd1 vccd1 vccd1 _12651_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _10470_/Y _09179_/C _11603_/S vssd1 vssd1 vccd1 vccd1 _11602_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12582_ _12993_/CLK _12582_/D vssd1 vssd1 vccd1 vccd1 _12582_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _12822_/Q _09180_/D _11533_/S vssd1 vssd1 vccd1 vccd1 _11533_/X sky130_fd_sc_hd__mux2_1
XPHY_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11464_ _12907_/Q _09243_/A _11469_/S vssd1 vssd1 vccd1 vccd1 _11464_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13203_ _13205_/CLK _13203_/D _06747_/X vssd1 vssd1 vccd1 vccd1 _13203_/Q sky130_fd_sc_hd__dfrtp_1
X_10415_ _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10418_/B sky130_fd_sc_hd__or2_1
XFILLER_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11395_ _10607_/Y _12410_/D _11404_/S vssd1 vssd1 vccd1 vccd1 _11395_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13134_ _12168_/X _13134_/D _07142_/X vssd1 vssd1 vccd1 vccd1 _13134_/Q sky130_fd_sc_hd__dfrtp_4
X_10346_ _10346_/A _10346_/B _10346_/C vssd1 vssd1 vccd1 vccd1 _10352_/C sky130_fd_sc_hd__or3_4
XFILLER_3_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13065_ _12165_/X _13065_/D _07343_/X vssd1 vssd1 vccd1 vccd1 _13065_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10277_ _10277_/A vssd1 vssd1 vccd1 vccd1 _10277_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_140_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12016_ _11097_/X _11092_/X _12200_/S vssd1 vssd1 vccd1 vccd1 _12016_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12918_ _12166_/X _12918_/D _07906_/X vssd1 vssd1 vccd1 vccd1 _12918_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_185_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12849_ _12849_/CLK _12849_/D _08094_/X vssd1 vssd1 vccd1 vccd1 _12849_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_181_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06370_ _06370_/A vssd1 vssd1 vccd1 vccd1 _06370_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08040_ _08040_/A vssd1 vssd1 vccd1 vccd1 _08040_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09991_ _09991_/A vssd1 vssd1 vccd1 vccd1 _09991_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_170_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08942_ _12426_/Q _12425_/Q vssd1 vssd1 vccd1 vccd1 _11370_/S sky130_fd_sc_hd__nor2_1
XFILLER_97_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08873_ _08882_/A vssd1 vssd1 vccd1 vccd1 _08873_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07824_ _12918_/Q vssd1 vssd1 vccd1 vccd1 _07824_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07755_ _12581_/Q _07755_/B vssd1 vssd1 vccd1 vccd1 _07756_/B sky130_fd_sc_hd__or2_1
XFILLER_84_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06706_ _06630_/X _06694_/X _06704_/X _06646_/X _06705_/Y vssd1 vssd1 vccd1 vccd1
+ _06707_/A sky130_fd_sc_hd__a32o_1
X_07686_ _07686_/A _07686_/B vssd1 vssd1 vccd1 vccd1 _07686_/X sky130_fd_sc_hd__or2_1
XFILLER_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09425_ _12465_/Q _10579_/A _09355_/Y _12415_/D vssd1 vssd1 vccd1 vccd1 _09425_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06637_ _12087_/X vssd1 vssd1 vccd1 vccd1 _06637_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _12396_/Q vssd1 vssd1 vccd1 vccd1 _09356_/Y sky130_fd_sc_hd__inv_2
X_06568_ _12178_/X _12177_/X _06562_/X _06563_/X _06567_/X vssd1 vssd1 vccd1 vccd1
+ _06569_/A sky130_fd_sc_hd__o32a_1
XFILLER_139_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_139_wb_clk_i _13253_/CLK vssd1 vssd1 vccd1 vccd1 _12886_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_100_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08307_ _12824_/Q _11599_/X _08307_/S vssd1 vssd1 vccd1 vccd1 _12824_/D sky130_fd_sc_hd__mux2_1
X_09287_ _09288_/A _09288_/B _10015_/B _09274_/B _09271_/X vssd1 vssd1 vccd1 vccd1
+ _12301_/D sky130_fd_sc_hd__a41o_1
XFILLER_166_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06499_ _12041_/X _06484_/X _12041_/X _06484_/X vssd1 vssd1 vccd1 vccd1 _06500_/B
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08238_ _08238_/A _08238_/B _08238_/C _08237_/X vssd1 vssd1 vccd1 vccd1 _08247_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_5_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08169_ _12820_/Q vssd1 vssd1 vccd1 vccd1 _10455_/B sky130_fd_sc_hd__inv_2
XFILLER_10_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10200_ _12885_/Q vssd1 vssd1 vccd1 vccd1 _10200_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11180_ vssd1 vssd1 vccd1 vccd1 _11180_/HI _11180_/LO sky130_fd_sc_hd__conb_1
X_10131_ _11969_/S _10527_/C _09982_/D _13078_/Q _10130_/X vssd1 vssd1 vccd1 vccd1
+ _10131_/X sky130_fd_sc_hd__a41o_1
XFILLER_121_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10062_ _10061_/Y _10028_/X _09890_/Y _10134_/A vssd1 vssd1 vccd1 vccd1 _10068_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10964_ _10962_/Y _10963_/Y _12536_/Q _12348_/Q vssd1 vssd1 vccd1 vccd1 _10976_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12703_ _12707_/CLK _12703_/D _08695_/X vssd1 vssd1 vccd1 vccd1 _12703_/Q sky130_fd_sc_hd__dfrtp_1
X_10895_ _10895_/A vssd1 vssd1 vccd1 vccd1 _10895_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ _13158_/CLK _12634_/D _08886_/X vssd1 vssd1 vccd1 vccd1 _12634_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12565_ _12570_/CLK _12565_/D vssd1 vssd1 vccd1 vccd1 _12565_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11516_ _12805_/Q _09185_/D _11546_/S vssd1 vssd1 vccd1 vccd1 _11516_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12496_ _12992_/CLK _12496_/D vssd1 vssd1 vccd1 vccd1 _12496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11447_ _12922_/Q _10794_/A _11449_/S vssd1 vssd1 vccd1 vccd1 _11447_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11378_ _10592_/X _12405_/D _11404_/S vssd1 vssd1 vccd1 vccd1 _11378_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10329_ _10331_/B vssd1 vssd1 vccd1 vccd1 _10329_/Y sky130_fd_sc_hd__inv_2
X_13117_ _12168_/X _13117_/D _07186_/X vssd1 vssd1 vccd1 vccd1 _13117_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13048_ _12165_/X _13048_/D _07387_/X vssd1 vssd1 vccd1 vccd1 _13048_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_67_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07540_ _12998_/Q _07531_/X _09186_/A _07532_/X _07538_/X vssd1 vssd1 vccd1 vccd1
+ _12998_/D sky130_fd_sc_hd__o221a_1
XFILLER_81_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07471_ _07473_/A vssd1 vssd1 vccd1 vccd1 _07471_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_50_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09210_ _12479_/Q _09207_/X _09243_/C _09208_/X vssd1 vssd1 vccd1 vccd1 _12479_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06422_ _12768_/Q vssd1 vssd1 vccd1 vccd1 _10714_/B sky130_fd_sc_hd__inv_2
XFILLER_34_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09141_ _12502_/Q _09141_/B vssd1 vssd1 vccd1 vccd1 _09142_/B sky130_fd_sc_hd__or2_1
XFILLER_33_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06353_ _06370_/A vssd1 vssd1 vccd1 vccd1 _06353_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_72_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09072_ _09072_/A _09072_/B _09072_/C vssd1 vssd1 vccd1 vccd1 _11030_/B sky130_fd_sc_hd__or3_4
X_06284_ _06269_/X _06281_/X _06283_/Y _13268_/Q _06273_/X vssd1 vssd1 vccd1 vccd1
+ _13268_/D sky130_fd_sc_hd__a32o_1
XFILLER_163_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08023_ _08025_/A vssd1 vssd1 vccd1 vccd1 _08040_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_200_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09974_ _09981_/A _10090_/A vssd1 vssd1 vccd1 vccd1 _10141_/A sky130_fd_sc_hd__or2_4
XFILLER_170_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08925_ _08925_/A _08925_/B vssd1 vssd1 vccd1 vccd1 _08926_/B sky130_fd_sc_hd__or2_1
XFILLER_103_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08856_ _08866_/A vssd1 vssd1 vccd1 vccd1 _08856_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_85_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07807_ _12899_/Q vssd1 vssd1 vccd1 vccd1 _10333_/A sky130_fd_sc_hd__clkinv_4
X_08787_ _12672_/Q vssd1 vssd1 vccd1 vccd1 _08787_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07738_ _12944_/Q _07729_/X _07737_/X vssd1 vssd1 vccd1 vccd1 _12944_/D sky130_fd_sc_hd__o21a_1
XFILLER_198_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07669_ _12952_/Q _12949_/Q _07658_/A vssd1 vssd1 vccd1 vccd1 _07669_/X sky130_fd_sc_hd__a21bo_1
XFILLER_41_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09408_ _12403_/D vssd1 vssd1 vccd1 vccd1 _09418_/A sky130_fd_sc_hd__inv_2
XFILLER_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ _12445_/Q vssd1 vssd1 vccd1 vccd1 _10680_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09339_ _12459_/Q _09337_/Y _09338_/Y _12409_/Q vssd1 vssd1 vccd1 vccd1 _09339_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ _12353_/CLK _12350_/D vssd1 vssd1 vccd1 vccd1 _12350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11301_ vssd1 vssd1 vccd1 vccd1 _11301_/HI _11301_/LO sky130_fd_sc_hd__conb_1
X_12281_ _10309_/X _12907_/Q _11877_/X _10307_/Y _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12297_/D sky130_fd_sc_hd__mux4_2
XFILLER_101_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11232_ vssd1 vssd1 vccd1 vccd1 _11232_/HI _11232_/LO sky130_fd_sc_hd__conb_1
XFILLER_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ vssd1 vssd1 vccd1 vccd1 _11163_/HI _11163_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_wb_clk_i clkbuf_4_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12376_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10114_ _10112_/Y _10090_/X _08445_/Y _10113_/X vssd1 vssd1 vccd1 vccd1 _10114_/X
+ sky130_fd_sc_hd__o22a_1
X_11094_ _06365_/X _11045_/A _08535_/A _10736_/X _07030_/X vssd1 vssd1 vccd1 vccd1
+ _11094_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput320 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 _07102_/A sky130_fd_sc_hd__clkbuf_1
Xinput331 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 _07990_/A sky130_fd_sc_hd__buf_2
Xinput342 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 input342/X sky130_fd_sc_hd__clkbuf_2
X_10045_ _10045_/A vssd1 vssd1 vccd1 vccd1 _10796_/A sky130_fd_sc_hd__buf_2
Xinput353 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 _10793_/A sky130_fd_sc_hd__buf_4
Xinput364 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _09293_/D sky130_fd_sc_hd__buf_1
XFILLER_64_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11996_ _11103_/X _11095_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _11996_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10947_ _10947_/A _10947_/B _10947_/C vssd1 vssd1 vccd1 vccd1 _10947_/Y sky130_fd_sc_hd__nor3_2
XFILLER_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10878_ _10877_/A _10876_/Y _10890_/B _10876_/A vssd1 vssd1 vccd1 vccd1 _12335_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _12769_/CLK _12617_/D _08960_/X vssd1 vssd1 vccd1 vccd1 _12617_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12548_ _12550_/CLK _12548_/D _09070_/X vssd1 vssd1 vccd1 vccd1 _12548_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_200_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12479_ _12480_/CLK _12479_/D vssd1 vssd1 vccd1 vccd1 _12479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06971_ _06971_/A _06971_/B vssd1 vssd1 vccd1 vccd1 _06971_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08710_ _08714_/A vssd1 vssd1 vccd1 vccd1 _08710_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09690_ _09690_/A vssd1 vssd1 vccd1 vccd1 _09690_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08641_ _11934_/X _08639_/X _12725_/Q _08640_/X vssd1 vssd1 vccd1 vccd1 _12725_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08572_ _12613_/Q _12614_/Q _09491_/A vssd1 vssd1 vccd1 vccd1 _09469_/A sky130_fd_sc_hd__or3_4
XFILLER_70_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07523_ _13004_/Q _07520_/Y _09226_/A _07520_/A _07522_/Y vssd1 vssd1 vccd1 vccd1
+ _13004_/D sky130_fd_sc_hd__o221a_1
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07454_ _07458_/A vssd1 vssd1 vccd1 vccd1 _07454_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_179_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06405_ _06403_/X _12208_/X _06396_/X _06404_/X vssd1 vssd1 vccd1 vccd1 _13241_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07385_ _07385_/A vssd1 vssd1 vccd1 vccd1 _07385_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_176_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06336_ _06336_/A vssd1 vssd1 vccd1 vccd1 _06336_/Y sky130_fd_sc_hd__clkinv_4
X_09124_ _09124_/A vssd1 vssd1 vccd1 vccd1 _09124_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09055_ _09058_/A _12151_/X vssd1 vssd1 vccd1 vccd1 _12562_/D sky130_fd_sc_hd__nor2b_1
XFILLER_175_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06267_ _06280_/A vssd1 vssd1 vccd1 vccd1 _06267_/X sky130_fd_sc_hd__clkbuf_1
X_08006_ _12883_/Q _07996_/X _08005_/X _07998_/X vssd1 vssd1 vccd1 vccd1 _12883_/D
+ sky130_fd_sc_hd__a22o_1
X_06198_ _06144_/A _06197_/B _06196_/X _06151_/B _06197_/X vssd1 vssd1 vccd1 vccd1
+ _06198_/X sky130_fd_sc_hd__o311a_1
XFILLER_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09957_ _08759_/Y _09952_/X _06212_/X _09949_/X _09950_/X vssd1 vssd1 vccd1 vccd1
+ _09957_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_106_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08908_ _12612_/Q vssd1 vssd1 vccd1 vccd1 _08908_/X sky130_fd_sc_hd__buf_2
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09888_ _12877_/Q _09478_/X _09475_/X vssd1 vssd1 vccd1 vccd1 _09888_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_46_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08839_ _08839_/A vssd1 vssd1 vccd1 vccd1 _08851_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _09961_/Y _12860_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11850_/X sky130_fd_sc_hd__mux2_1
XPHY_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_154_wb_clk_i clkbuf_4_8_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12357_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10801_ _12511_/Q _12323_/Q _12511_/Q _12323_/Q vssd1 vssd1 vccd1 vccd1 _10801_/X
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _12136_/X _11780_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11781_/X sky130_fd_sc_hd__mux2_1
XPHY_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10732_ _11111_/A vssd1 vssd1 vccd1 vccd1 _10732_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10663_ _12426_/Q _12425_/Q _12427_/Q vssd1 vssd1 vccd1 vccd1 _10663_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12402_ _12415_/CLK _12402_/D vssd1 vssd1 vccd1 vccd1 _12402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10594_ _10594_/A _10594_/B vssd1 vssd1 vccd1 vccd1 _10594_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12333_ _12535_/CLK _12333_/D vssd1 vssd1 vccd1 vccd1 _12333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12264_ _12263_/X _12652_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12264_/X sky130_fd_sc_hd__mux2_2
XFILLER_107_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11215_ vssd1 vssd1 vccd1 vccd1 _11215_/HI _11215_/LO sky130_fd_sc_hd__conb_1
X_12195_ _10757_/Y _06491_/A _12764_/Q vssd1 vssd1 vccd1 vccd1 _12195_/X sky130_fd_sc_hd__mux2_2
X_11146_ _11146_/A vssd1 vssd1 vccd1 vccd1 _11146_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11077_ _11077_/A vssd1 vssd1 vccd1 vccd1 _11077_/X sky130_fd_sc_hd__clkbuf_2
Xinput150 la_data_in[85] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_hd__buf_1
Xinput161 la_data_in[95] vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_hd__buf_1
Xinput172 la_oenb[104] vssd1 vssd1 vccd1 vccd1 input172/X sky130_fd_sc_hd__buf_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10028_ _10137_/A vssd1 vssd1 vccd1 vccd1 _10028_/X sky130_fd_sc_hd__clkbuf_2
Xinput183 la_oenb[114] vssd1 vssd1 vccd1 vccd1 input183/X sky130_fd_sc_hd__buf_1
Xinput194 la_oenb[124] vssd1 vssd1 vccd1 vccd1 input194/X sky130_fd_sc_hd__buf_1
XFILLER_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11979_ _10189_/Y _12795_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11979_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07170_ _07253_/A vssd1 vssd1 vccd1 vccd1 _07183_/A sky130_fd_sc_hd__buf_2
XFILLER_191_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06121_ _12718_/Q _12686_/Q _12944_/Q _06120_/X vssd1 vssd1 vccd1 vccd1 _06122_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06052_ _12738_/Q _12706_/Q _12738_/Q _12706_/Q vssd1 vssd1 vccd1 vccd1 _06056_/A
+ sky130_fd_sc_hd__a2bb2oi_2
Xoutput602 _12288_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_154_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09811_ _13225_/Q _13224_/Q _06529_/Y _06533_/Y vssd1 vssd1 vccd1 vccd1 _09812_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_114_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09742_ _09742_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__or2_1
X_06954_ _10759_/A _06954_/B vssd1 vssd1 vccd1 vccd1 _06954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09673_ _09673_/A _09673_/B vssd1 vssd1 vccd1 vccd1 _09714_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06885_ _06916_/A vssd1 vssd1 vccd1 vccd1 _06885_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_94_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08624_ _08685_/A vssd1 vssd1 vccd1 vccd1 _08624_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _12610_/Q vssd1 vssd1 vccd1 vccd1 _08740_/A sky130_fd_sc_hd__inv_2
XFILLER_36_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07506_ _07609_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _13007_/D sky130_fd_sc_hd__nor2_1
XFILLER_39_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08486_ _13059_/Q _12910_/Q _13059_/Q _12910_/Q vssd1 vssd1 vccd1 vccd1 _08486_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07437_ _07443_/A vssd1 vssd1 vccd1 vccd1 _07437_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12960_/CLK
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07368_ _07368_/A vssd1 vssd1 vccd1 vccd1 _07368_/X sky130_fd_sc_hd__buf_2
XFILLER_182_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09107_ _09115_/A vssd1 vssd1 vccd1 vccd1 _09107_/X sky130_fd_sc_hd__clkbuf_2
X_06319_ _06344_/A vssd1 vssd1 vccd1 vccd1 _06319_/X sky130_fd_sc_hd__clkbuf_1
X_07299_ _09186_/B vssd1 vssd1 vccd1 vccd1 _07562_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09038_ _13002_/Q vssd1 vssd1 vccd1 vccd1 _09038_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11000_ _11000_/A _11000_/B _11000_/C _11000_/D vssd1 vssd1 vccd1 vccd1 _11000_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_81_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ _12951_/CLK _12951_/D vssd1 vssd1 vccd1 vccd1 _12951_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11902_ _06491_/A _10757_/Y _12764_/Q vssd1 vssd1 vccd1 vccd1 _12201_/S sky130_fd_sc_hd__mux2_8
XPHY_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _12886_/CLK _12882_/D _08008_/X vssd1 vssd1 vccd1 vccd1 _12882_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_46_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11833_ _09933_/Y _12858_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11833_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _09184_/B _11763_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11764_/X sky130_fd_sc_hd__mux2_1
XPHY_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10715_ _12769_/Q _12768_/Q vssd1 vssd1 vccd1 vccd1 _10715_/Y sky130_fd_sc_hd__nor2_2
XFILLER_158_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _11402_/X _09179_/A _11703_/S vssd1 vssd1 vccd1 vccd1 _11695_/X sky130_fd_sc_hd__mux2_1
XPHY_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ _11905_/X _10649_/B vssd1 vssd1 vccd1 vccd1 _10646_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10577_ _10583_/A _11390_/X vssd1 vssd1 vccd1 vccd1 _10577_/Y sky130_fd_sc_hd__nor2b_1
Xclkbuf_leaf_51_wb_clk_i clkbuf_4_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13001_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ _12987_/CLK _12316_/D vssd1 vssd1 vccd1 vccd1 _12316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12247_ _12778_/Q _12851_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12247_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12178_ _11138_/X _11134_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _12178_/X sky130_fd_sc_hd__mux2_2
XFILLER_150_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11129_ _11129_/A vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06670_ _12048_/X _12047_/X _06664_/X _06665_/X _06669_/X vssd1 vssd1 vccd1 vccd1
+ _06671_/A sky130_fd_sc_hd__o32a_1
XFILLER_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08340_ _12810_/Q _11585_/X _08349_/S vssd1 vssd1 vccd1 vccd1 _12810_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08271_ _08271_/A _09969_/B _09296_/A vssd1 vssd1 vccd1 vccd1 _08271_/Y sky130_fd_sc_hd__nor3_4
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07222_ _11571_/X _07218_/X _13106_/Q _07219_/X vssd1 vssd1 vccd1 vccd1 _13106_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07153_ _11531_/X _07145_/X _13130_/Q _07146_/X vssd1 vssd1 vccd1 vccd1 _13130_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06104_ _12724_/Q _12692_/Q _12724_/Q _12692_/Q vssd1 vssd1 vccd1 vccd1 _06108_/A
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_118_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07084_ _13079_/Q vssd1 vssd1 vccd1 vccd1 _07084_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput410 _11192_/LO vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput421 _11202_/LO vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__clkbuf_2
Xoutput432 _11212_/LO vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06035_ _06035_/A _06035_/B vssd1 vssd1 vccd1 vccd1 _06035_/X sky130_fd_sc_hd__or2_1
Xoutput443 _11152_/HI vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput454 _11323_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__clkbuf_2
Xoutput465 _11333_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__clkbuf_2
Xoutput476 _11343_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__clkbuf_2
Xoutput487 _11237_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput498 _11247_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__clkbuf_2
X_07986_ _07986_/A vssd1 vssd1 vccd1 vccd1 _07986_/X sky130_fd_sc_hd__buf_2
XFILLER_41_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09725_ _09725_/A vssd1 vssd1 vccd1 vccd1 _09725_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06937_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06937_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_68_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09656_ _09655_/A _09655_/B _09671_/A vssd1 vssd1 vccd1 vccd1 _09657_/A sky130_fd_sc_hd__a21bo_1
X_06868_ _07026_/A vssd1 vssd1 vccd1 vccd1 _06916_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_1_wb_clk_i clkbuf_2_3_1_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_1
X_08607_ _08715_/A vssd1 vssd1 vccd1 vccd1 _08685_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09587_ _13184_/Q vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__inv_2
X_06799_ _06797_/X _06798_/X _06797_/X _06798_/X vssd1 vssd1 vccd1 vccd1 _06804_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08642_/A vssd1 vssd1 vccd1 vccd1 _08569_/A sky130_fd_sc_hd__buf_4
XPHY_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _08461_/Y _10318_/A _13067_/Q _07824_/Y vssd1 vssd1 vccd1 vccd1 _08473_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10500_ _12505_/Q _09144_/B _09145_/B vssd1 vssd1 vccd1 vccd1 _10500_/X sky130_fd_sc_hd__a21bo_1
XPHY_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11480_ _12923_/Q _10793_/B _11481_/S vssd1 vssd1 vccd1 vccd1 _11480_/X sky130_fd_sc_hd__mux2_1
XPHY_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10431_ _10431_/A _10431_/B _10474_/A vssd1 vssd1 vccd1 vccd1 _10431_/Y sky130_fd_sc_hd__nor3_2
XFILLER_195_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13150_ _13152_/CLK _13150_/D _07073_/X vssd1 vssd1 vccd1 vccd1 _13150_/Q sky130_fd_sc_hd__dfrtp_2
X_10362_ _10368_/A _10362_/B _10368_/D vssd1 vssd1 vccd1 vccd1 _10363_/A sky130_fd_sc_hd__or3_4
XFILLER_3_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12101_ _10667_/X _08949_/B _12101_/S vssd1 vssd1 vccd1 vccd1 _12101_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13081_ _13081_/CLK _13081_/D _07283_/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfrtp_2
X_10293_ _13095_/Q _10276_/X _13127_/Q _10277_/X vssd1 vssd1 vccd1 vccd1 _10293_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12032_ _06698_/B _11102_/X _12185_/S vssd1 vssd1 vccd1 vccd1 _12032_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12934_ _12973_/CLK _12934_/D vssd1 vssd1 vccd1 vccd1 _12934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12865_ _12868_/CLK _12865_/D _08051_/X vssd1 vssd1 vccd1 vccd1 _12865_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _12096_/X _12492_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11816_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12864_/CLK _12796_/D _08377_/X vssd1 vssd1 vccd1 vccd1 _12796_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_109_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11747_ _11374_/X _12471_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11747_/X sky130_fd_sc_hd__mux2_1
XPHY_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11678_ _11677_/X _11382_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12381_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10629_ _11890_/X vssd1 vssd1 vccd1 vccd1 _10629_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13279_ _13279_/CLK _13279_/D _06221_/X vssd1 vssd1 vccd1 vccd1 _13279_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07840_ _13021_/Q _07839_/X _13021_/Q _07839_/X vssd1 vssd1 vccd1 vccd1 _07840_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_151_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07771_ _12937_/Q _11648_/S _12938_/Q _07769_/X _07569_/X vssd1 vssd1 vccd1 vccd1
+ _12938_/D sky130_fd_sc_hd__a221o_1
XFILLER_83_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09510_ _13151_/Q vssd1 vssd1 vccd1 vccd1 _09510_/Y sky130_fd_sc_hd__inv_2
X_06722_ _06750_/A vssd1 vssd1 vccd1 vccd1 _06722_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _09441_/A _10527_/B _10527_/C vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__and3_2
X_06653_ _06640_/X _06644_/X _06645_/X vssd1 vssd1 vccd1 vccd1 _06653_/X sky130_fd_sc_hd__a21bo_1
XFILLER_91_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09372_ _09349_/Y _12413_/Q _09362_/Y _12398_/Q vssd1 vssd1 vccd1 vccd1 _09372_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06584_ _10745_/A vssd1 vssd1 vccd1 vccd1 _07007_/A sky130_fd_sc_hd__inv_2
XFILLER_36_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08323_ _08353_/S vssd1 vssd1 vccd1 vccd1 _08335_/S sky130_fd_sc_hd__buf_2
XFILLER_123_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08254_ _12842_/Q _08251_/X _07290_/X _11417_/S vssd1 vssd1 vccd1 vccd1 _12842_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07205_ _11578_/X _07201_/X _13113_/Q _07204_/X vssd1 vssd1 vccd1 vccd1 _13113_/D
+ sky130_fd_sc_hd__a22o_1
X_08185_ _08107_/Y _10484_/A _08183_/Y _12826_/Q _08184_/X vssd1 vssd1 vccd1 vccd1
+ _08190_/C sky130_fd_sc_hd__o221a_1
XFILLER_192_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07136_ _11538_/X _07130_/X _13137_/Q _07131_/X vssd1 vssd1 vccd1 vccd1 _13137_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07067_ _07053_/X _07058_/X _06323_/Y _13153_/Q _07059_/X vssd1 vssd1 vccd1 vccd1
+ _13153_/D sky130_fd_sc_hd__a32o_1
XFILLER_161_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06018_ _12548_/Q _09282_/A _11031_/A vssd1 vssd1 vccd1 vccd1 _08562_/B sky130_fd_sc_hd__o21ai_4
XFILLER_133_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07969_ _09986_/D vssd1 vssd1 vccd1 vccd1 _09982_/D sky130_fd_sc_hd__buf_2
XFILLER_101_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09708_ _09708_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _09709_/A sky130_fd_sc_hd__or2_1
XFILLER_28_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10980_ _10980_/A _10980_/B vssd1 vssd1 vccd1 vccd1 _10980_/Y sky130_fd_sc_hd__nand2_2
XFILLER_28_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09639_ _13194_/Q _09638_/A _09637_/Y _09638_/Y vssd1 vssd1 vccd1 vccd1 _09640_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ _12653_/CLK _12650_/D _08844_/X vssd1 vssd1 vccd1 vccd1 _12650_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _10466_/X _09179_/D _11603_/S vssd1 vssd1 vccd1 vccd1 _11601_/X sky130_fd_sc_hd__mux2_1
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12581_ _12993_/CLK _12581_/D vssd1 vssd1 vccd1 vccd1 _12581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11532_ _12821_/Q _09179_/A _11533_/S vssd1 vssd1 vccd1 vccd1 _11532_/X sky130_fd_sc_hd__mux2_1
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11463_ _12906_/Q input333/X _11469_/S vssd1 vssd1 vccd1 vccd1 _11463_/X sky130_fd_sc_hd__mux2_1
XPHY_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13202_ _13205_/CLK _13202_/D _06750_/X vssd1 vssd1 vccd1 vccd1 _13202_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_139_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10414_ _08113_/X _10413_/B _10415_/B _10407_/X vssd1 vssd1 vccd1 vccd1 _10414_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11394_ _11048_/X _11044_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _11394_/X sky130_fd_sc_hd__mux2_1
X_13133_ _12168_/X _13133_/D _07144_/X vssd1 vssd1 vccd1 vccd1 _13133_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10345_ _12903_/Q _10344_/B _10346_/B _10346_/C _10320_/X vssd1 vssd1 vccd1 vccd1
+ _10345_/X sky130_fd_sc_hd__o221a_1
XFILLER_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13064_ _12165_/X _13064_/D _07345_/X vssd1 vssd1 vccd1 vccd1 _13064_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10276_ _10276_/A vssd1 vssd1 vccd1 vccd1 _10276_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12015_ _11081_/X _11073_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12015_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12917_ _12166_/X _12917_/D _07909_/X vssd1 vssd1 vccd1 vccd1 _12917_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12848_ _12849_/CLK _12848_/D _08096_/X vssd1 vssd1 vccd1 vccd1 _12848_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12779_ _12779_/CLK _12779_/D _08423_/X vssd1 vssd1 vccd1 vccd1 _12779_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09990_ _10001_/A vssd1 vssd1 vccd1 vccd1 _09991_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08941_ _12428_/Q vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__inv_2
XFILLER_170_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08872_ _07747_/X _06346_/Y _08837_/A _12639_/Q vssd1 vssd1 vccd1 vccd1 _12639_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07823_ _12895_/Q vssd1 vssd1 vccd1 vccd1 _07823_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07754_ _12580_/Q _12579_/Q vssd1 vssd1 vccd1 vccd1 _07755_/B sky130_fd_sc_hd__or2_1
XFILLER_38_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06705_ _13208_/Q vssd1 vssd1 vccd1 vccd1 _06705_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07685_ _07685_/A _07685_/B _07685_/C _07685_/D vssd1 vssd1 vccd1 vccd1 _07686_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09424_ _12401_/D vssd1 vssd1 vccd1 vccd1 _10579_/A sky130_fd_sc_hd__inv_2
XFILLER_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06636_ _06636_/A vssd1 vssd1 vccd1 vccd1 _11071_/A sky130_fd_sc_hd__clkbuf_2
X_09355_ _12546_/Q vssd1 vssd1 vccd1 vccd1 _09355_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06567_ _06564_/X _06565_/X _12170_/X _06566_/X vssd1 vssd1 vccd1 vccd1 _06567_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_138_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08306_ _08311_/A vssd1 vssd1 vccd1 vccd1 _08306_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_139_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09286_ _09286_/A _09286_/B vssd1 vssd1 vccd1 vccd1 _12300_/D sky130_fd_sc_hd__nand2_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06498_ _12040_/X _06494_/Y _06495_/Y _06497_/Y vssd1 vssd1 vccd1 vccd1 _06500_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_166_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08237_ _08233_/X _08237_/B _08237_/C _08237_/D vssd1 vssd1 vccd1 vccd1 _08237_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_119_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08168_ _13143_/Q _10482_/A _13138_/Q _08164_/Y vssd1 vssd1 vccd1 vccd1 _08175_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_108_wb_clk_i _12726_/CLK vssd1 vssd1 vccd1 vccd1 _12735_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_146_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07119_ _11545_/X _07113_/X _13144_/Q _07116_/X vssd1 vssd1 vccd1 vccd1 _13144_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08099_ _12847_/Q _08082_/A _07304_/X _08083_/A vssd1 vssd1 vccd1 vccd1 _12847_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10130_ _13086_/Q _10276_/A _13118_/Q _10277_/A vssd1 vssd1 vccd1 vccd1 _10130_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10061_ _12846_/Q vssd1 vssd1 vccd1 vccd1 _10061_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10963_ _12348_/Q vssd1 vssd1 vccd1 vccd1 _10963_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12702_ _12716_/CLK _12702_/D _08697_/X vssd1 vssd1 vccd1 vccd1 _12702_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10894_ _12526_/Q _12338_/Q _12526_/Q _12338_/Q vssd1 vssd1 vccd1 vccd1 _10921_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12633_ _13158_/CLK _12633_/D _08888_/X vssd1 vssd1 vccd1 vccd1 _12633_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12564_ _12570_/CLK _12564_/D vssd1 vssd1 vccd1 vccd1 _12564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11515_ _12804_/Q _09184_/A _11546_/S vssd1 vssd1 vccd1 vccd1 _11515_/X sky130_fd_sc_hd__mux2_1
XPHY_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12495_ _12986_/CLK _12495_/D vssd1 vssd1 vccd1 vccd1 _12495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11446_ _12921_/Q _10794_/B _11449_/S vssd1 vssd1 vccd1 vccd1 _11446_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11377_ _10594_/Y _12406_/D _11404_/S vssd1 vssd1 vccd1 vccd1 _11377_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13116_ _12168_/X _13116_/D _07188_/X vssd1 vssd1 vccd1 vccd1 _13116_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10328_ _10328_/A _10328_/B vssd1 vssd1 vccd1 vccd1 _10331_/B sky130_fd_sc_hd__or2_1
XFILLER_112_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13047_ _12165_/X _13047_/D _07389_/X vssd1 vssd1 vccd1 vccd1 _13047_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10259_ _09925_/Y _09968_/X _10250_/X _10258_/X vssd1 vssd1 vccd1 vccd1 _10259_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_65_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07470_ _11459_/X _07459_/X _13018_/Q _07460_/X vssd1 vssd1 vccd1 vccd1 _13018_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06421_ _12769_/Q vssd1 vssd1 vccd1 vccd1 _10714_/A sky130_fd_sc_hd__inv_2
XFILLER_201_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09140_ _12501_/Q _09140_/B vssd1 vssd1 vccd1 vccd1 _09141_/B sky130_fd_sc_hd__or2_1
X_06352_ _07742_/B _06281_/A _06351_/X _13255_/Q _06306_/A vssd1 vssd1 vccd1 vccd1
+ _13255_/D sky130_fd_sc_hd__a32o_1
XFILLER_33_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_wb_clk_i _12844_/CLK vssd1 vssd1 vccd1 vccd1 _12864_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_187_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09071_ _09071_/A _09071_/B _09071_/C _09071_/D vssd1 vssd1 vccd1 vccd1 _09072_/B
+ sky130_fd_sc_hd__or4_4
X_06283_ _06283_/A vssd1 vssd1 vccd1 vccd1 _06283_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_163_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08022_ _10090_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08025_/A sky130_fd_sc_hd__or2_1
XFILLER_116_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09973_ _12876_/Q vssd1 vssd1 vccd1 vccd1 _09973_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08924_ _12417_/Q vssd1 vssd1 vccd1 vccd1 _08925_/B sky130_fd_sc_hd__inv_2
XFILLER_130_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08855_ _08963_/A vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07806_ _07799_/Y _07800_/X _07801_/Y _10388_/A _07805_/X vssd1 vssd1 vccd1 vccd1
+ _07819_/B sky130_fd_sc_hd__a221o_1
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08786_ _08789_/A vssd1 vssd1 vccd1 vccd1 _08786_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_84_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07737_ _07737_/A vssd1 vssd1 vccd1 vccd1 _07737_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07668_ _07684_/A _07668_/B _07668_/C _07685_/D vssd1 vssd1 vccd1 vccd1 _07672_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_168_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09407_ _12544_/Q _10619_/A _12457_/Q _10603_/A _09406_/X vssd1 vssd1 vccd1 vccd1
+ _09431_/A sky130_fd_sc_hd__a221o_1
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06619_ _06625_/A _06625_/B vssd1 vssd1 vccd1 vccd1 _06620_/B sky130_fd_sc_hd__and2_1
XFILLER_186_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07599_ _12601_/Q vssd1 vssd1 vccd1 vccd1 _07599_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09338_ _12457_/Q vssd1 vssd1 vccd1 vccd1 _09338_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09269_ _09269_/A _12302_/Q _09271_/C vssd1 vssd1 vccd1 vccd1 _09269_/X sky130_fd_sc_hd__and3_1
XFILLER_194_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11300_ vssd1 vssd1 vccd1 vccd1 _11300_/HI _11300_/LO sky130_fd_sc_hd__conb_1
XFILLER_126_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12280_ _10294_/X _12906_/Q _11876_/X _10292_/Y _12282_/S0 _11348_/S vssd1 vssd1
+ vccd1 vccd1 _12296_/D sky130_fd_sc_hd__mux4_2
XFILLER_193_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11231_ vssd1 vssd1 vccd1 vccd1 _11231_/HI _11231_/LO sky130_fd_sc_hd__conb_1
XFILLER_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11162_ vssd1 vssd1 vccd1 vccd1 _11162_/HI _11162_/LO sky130_fd_sc_hd__conb_1
XFILLER_171_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10113_ _10113_/A vssd1 vssd1 vccd1 vccd1 _10113_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11093_ _11033_/X _11077_/X _06397_/X _11086_/X _11087_/X vssd1 vssd1 vccd1 vccd1
+ _11093_/X sky130_fd_sc_hd__a221o_1
XFILLER_150_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput310 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 _07097_/D sky130_fd_sc_hd__clkbuf_1
Xinput321 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _11969_/S sky130_fd_sc_hd__buf_6
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput332 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 _07986_/A sky130_fd_sc_hd__clkbuf_4
X_10044_ _10090_/A vssd1 vssd1 vccd1 vccd1 _10045_/A sky130_fd_sc_hd__buf_2
Xinput343 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 _09179_/D sky130_fd_sc_hd__buf_6
XFILLER_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_76_wb_clk_i _13219_/CLK vssd1 vssd1 vccd1 vccd1 _13201_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput354 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 input354/X sky130_fd_sc_hd__buf_1
XFILLER_48_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput365 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _07094_/A sky130_fd_sc_hd__buf_1
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11995_ _11059_/X _11053_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _11995_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10946_ _12531_/Q _12343_/Q _12530_/Q _12342_/Q vssd1 vssd1 vccd1 vccd1 _10946_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10877_ _10877_/A vssd1 vssd1 vccd1 vccd1 _10890_/B sky130_fd_sc_hd__inv_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ _12888_/CLK _12616_/D _08961_/X vssd1 vssd1 vccd1 vccd1 _12616_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12547_ _12547_/CLK _12547_/D vssd1 vssd1 vccd1 vccd1 _12547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12478_ _12480_/CLK _12478_/D vssd1 vssd1 vccd1 vccd1 _12478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11429_ _12904_/Q _09244_/B _11433_/S vssd1 vssd1 vccd1 vccd1 _11429_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06970_ _06977_/A _06977_/B vssd1 vssd1 vccd1 vccd1 _06971_/B sky130_fd_sc_hd__and2_1
XFILLER_101_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08640_ _08686_/A vssd1 vssd1 vccd1 vccd1 _08640_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08571_ _12611_/Q _09547_/A vssd1 vssd1 vccd1 vccd1 _09491_/A sky130_fd_sc_hd__or2_4
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _07522_/A _07522_/B vssd1 vssd1 vccd1 vccd1 _07522_/Y sky130_fd_sc_hd__nor2_2
XFILLER_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07453_ _11466_/X _07444_/X _13025_/Q _07445_/X vssd1 vssd1 vccd1 vccd1 _13025_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06404_ _13241_/Q vssd1 vssd1 vccd1 vccd1 _06404_/X sky130_fd_sc_hd__buf_2
XFILLER_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07384_ _07384_/A vssd1 vssd1 vccd1 vccd1 _07384_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09123_ _09123_/A vssd1 vssd1 vccd1 vccd1 _09123_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06335_ _06125_/C _06125_/B _06125_/C _06125_/B vssd1 vssd1 vccd1 vccd1 _06336_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_191_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09054_ _09058_/A _12152_/X vssd1 vssd1 vccd1 vccd1 _12563_/D sky130_fd_sc_hd__nor2b_1
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06266_ _06263_/Y _06247_/X _06217_/A _06265_/X vssd1 vssd1 vccd1 vccd1 _13271_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_159_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08005_ _09184_/B vssd1 vssd1 vccd1 vccd1 _08005_/X sky130_fd_sc_hd__buf_2
XFILLER_116_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06197_ _06197_/A _06197_/B vssd1 vssd1 vccd1 vccd1 _06197_/X sky130_fd_sc_hd__or2_1
XFILLER_144_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ _08763_/Y _09952_/X _06218_/X _09949_/X _09950_/X vssd1 vssd1 vccd1 vccd1
+ _09956_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_77_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08907_ _08912_/A vssd1 vssd1 vccd1 vccd1 _08907_/X sky130_fd_sc_hd__clkbuf_1
X_09887_ _11958_/S vssd1 vssd1 vccd1 vccd1 _11831_/S sky130_fd_sc_hd__buf_6
XFILLER_100_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08838_ _07746_/X _06271_/Y _12653_/Q _08837_/X vssd1 vssd1 vccd1 vccd1 _12653_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _08769_/A vssd1 vssd1 vccd1 vccd1 _08769_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10800_ _10799_/A _10799_/B _10799_/Y vssd1 vssd1 vccd1 vccd1 _12322_/D sky130_fd_sc_hd__a21oi_1
XPHY_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _09243_/C _11779_/X _11817_/S vssd1 vssd1 vccd1 vccd1 _11780_/X sky130_fd_sc_hd__mux2_1
XPHY_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ _10788_/A vssd1 vssd1 vccd1 vccd1 _10731_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10662_ _12426_/Q _12425_/Q vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__and2_1
XFILLER_90_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ _12464_/CLK _12401_/D vssd1 vssd1 vccd1 vccd1 _12401_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_123_wb_clk_i _12716_/CLK vssd1 vssd1 vccd1 vccd1 _12682_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10593_ _10525_/A _09390_/Y _09384_/Y _12403_/D _10586_/A vssd1 vssd1 vccd1 vccd1
+ _10594_/B sky130_fd_sc_hd__o32a_1
XFILLER_127_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12332_ _12535_/CLK _12332_/D vssd1 vssd1 vccd1 vccd1 _12332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ _12786_/Q _12859_/Q _12617_/Q vssd1 vssd1 vccd1 vccd1 _12263_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11214_ vssd1 vssd1 vccd1 vccd1 _11214_/HI _11214_/LO sky130_fd_sc_hd__conb_1
XFILLER_141_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12194_ _06451_/Y _10734_/X _12199_/S vssd1 vssd1 vccd1 vccd1 _12194_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11145_ _11145_/A vssd1 vssd1 vccd1 vccd1 _11145_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11076_ _11033_/X _11075_/X _06397_/X _10751_/X _10752_/X vssd1 vssd1 vccd1 vccd1
+ _11076_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput140 la_data_in[76] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_hd__buf_1
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput151 la_data_in[86] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_hd__buf_1
Xinput162 la_data_in[96] vssd1 vssd1 vccd1 vccd1 input162/X sky130_fd_sc_hd__buf_1
X_10027_ _12845_/Q vssd1 vssd1 vccd1 vccd1 _10027_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput173 la_oenb[105] vssd1 vssd1 vccd1 vccd1 input173/X sky130_fd_sc_hd__buf_1
Xinput184 la_oenb[115] vssd1 vssd1 vccd1 vccd1 input184/X sky130_fd_sc_hd__buf_1
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput195 la_oenb[125] vssd1 vssd1 vccd1 vccd1 input195/X sky130_fd_sc_hd__buf_1
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11978_ _10172_/Y _12794_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11978_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10929_ _12343_/Q vssd1 vssd1 vccd1 vccd1 _10930_/B sky130_fd_sc_hd__inv_2
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06120_ _12718_/Q _12686_/Q _12718_/Q _12686_/Q vssd1 vssd1 vccd1 vccd1 _06120_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_172_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06051_ _06051_/A _06050_/X vssd1 vssd1 vccd1 vccd1 _06209_/A sky130_fd_sc_hd__or2b_2
Xoutput603 _12289_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09810_ _13226_/Q vssd1 vssd1 vccd1 vccd1 _09810_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09741_ _13213_/Q _09740_/A _06659_/Y _09740_/Y vssd1 vssd1 vccd1 vccd1 _09742_/B
+ sky130_fd_sc_hd__a22o_2
X_06953_ _11077_/A vssd1 vssd1 vccd1 vccd1 _10759_/A sky130_fd_sc_hd__buf_2
XFILLER_189_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09672_ _09671_/A _09671_/B _09671_/Y vssd1 vssd1 vccd1 vccd1 _09713_/A sky130_fd_sc_hd__a21o_1
XFILLER_55_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06884_ _06829_/X _06870_/Y _06769_/X _06883_/Y vssd1 vssd1 vccd1 vccd1 _13189_/D
+ sky130_fd_sc_hd__o22ai_1
X_08623_ _08623_/A vssd1 vssd1 vccd1 vccd1 _08623_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08554_ _08556_/D _09259_/A vssd1 vssd1 vccd1 vccd1 _12616_/D sky130_fd_sc_hd__nor2_2
XPHY_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07505_ _07497_/Y _09227_/B _07522_/B _11982_/X _09284_/C vssd1 vssd1 vccd1 vccd1
+ _07506_/B sky130_fd_sc_hd__o32a_1
XFILLER_165_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08485_ _13056_/Q vssd1 vssd1 vccd1 vccd1 _08485_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07436_ _11473_/X _07429_/X _13032_/Q _07430_/X vssd1 vssd1 vccd1 vccd1 _13032_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07367_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07367_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_109_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09106_ _12530_/Q _09099_/X input341/X _09100_/X vssd1 vssd1 vccd1 vccd1 _12530_/D
+ sky130_fd_sc_hd__a22o_1
X_06318_ _06416_/A vssd1 vssd1 vccd1 vccd1 _06344_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07298_ _07302_/A vssd1 vssd1 vccd1 vccd1 _07298_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_108_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09037_ _12600_/Q _12572_/Q vssd1 vssd1 vccd1 vccd1 _09037_/X sky130_fd_sc_hd__or2_2
X_06249_ _06246_/Y _06247_/X _06217_/A _06248_/X vssd1 vssd1 vccd1 vccd1 _13274_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_191_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09939_ _12892_/Q _09939_/B vssd1 vssd1 vccd1 vccd1 _09950_/A sky130_fd_sc_hd__or2_2
X_12950_ _12955_/CLK _12950_/D vssd1 vssd1 vccd1 vccd1 _12950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11901_ _10762_/X _10764_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12881_ _12886_/CLK _12881_/D _08010_/X vssd1 vssd1 vccd1 vccd1 _12881_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _09930_/Y _12857_/Q _11851_/S vssd1 vssd1 vccd1 vccd1 _11832_/X sky130_fd_sc_hd__mux2_1
XPHY_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11763_ _12107_/X _12475_/Q _12142_/S vssd1 vssd1 vccd1 vccd1 _11763_/X sky130_fd_sc_hd__mux2_1
XPHY_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10714_/A _10714_/B vssd1 vssd1 vccd1 vccd1 _10714_/Y sky130_fd_sc_hd__nor2_1
XPHY_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _11693_/X _11405_/X _11704_/S vssd1 vssd1 vccd1 vccd1 _12389_/D sky130_fd_sc_hd__mux2_1
XPHY_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10645_ _11905_/X vssd1 vssd1 vccd1 vccd1 _10645_/Y sky130_fd_sc_hd__inv_2
XPHY_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10576_ _12399_/D _12400_/D _10579_/B vssd1 vssd1 vccd1 vccd1 _10576_/X sky130_fd_sc_hd__o21a_1
XFILLER_166_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12315_ _12987_/CLK _12315_/D vssd1 vssd1 vccd1 vccd1 _12315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12246_ _12245_/X _12643_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_91_wb_clk_i _13235_/CLK vssd1 vssd1 vccd1 vccd1 _13170_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12177_ _11137_/X _11133_/X _12202_/S vssd1 vssd1 vccd1 vccd1 _12177_/X sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_20_wb_clk_i _12468_/CLK vssd1 vssd1 vccd1 vccd1 _12492_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_111_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11128_ _13241_/Q _06425_/A _10696_/A _10717_/A _06430_/A vssd1 vssd1 vccd1 vccd1
+ _11129_/A sky130_fd_sc_hd__o221a_1
XFILLER_111_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11059_ _10779_/X _11037_/X _06389_/X _11058_/X _11038_/X vssd1 vssd1 vccd1 vccd1
+ _11059_/X sky130_fd_sc_hd__a221o_1
XFILLER_97_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08270_ _13078_/Q _08275_/A _08269_/Y vssd1 vssd1 vccd1 vccd1 _10411_/A sky130_fd_sc_hd__o21ai_4
XFILLER_60_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07221_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07221_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07152_ _07152_/A vssd1 vssd1 vccd1 vccd1 _07152_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06103_ _06103_/A _06103_/B vssd1 vssd1 vccd1 vccd1 _06130_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07083_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput400 _11345_/X vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__clkbuf_2
Xoutput411 _11193_/LO vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput422 _11203_/LO vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06034_ _06032_/Y _06033_/Y _12747_/Q _12715_/Q vssd1 vssd1 vccd1 vccd1 _06035_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput433 _11213_/LO vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput444 _12606_/Q vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__clkbuf_2
Xoutput455 _11324_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__clkbuf_2
Xoutput466 _11334_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__clkbuf_2
XFILLER_160_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput477 _11228_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput488 _11238_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput499 _11248_/LO vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__clkbuf_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07985_ _07985_/A vssd1 vssd1 vccd1 vccd1 _07985_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09724_ _13209_/Q vssd1 vssd1 vccd1 vccd1 _09724_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06936_ _06829_/X _09604_/B _06459_/X _06935_/Y vssd1 vssd1 vccd1 vccd1 _13183_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_28_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09655_ _09655_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__or2_2
X_06867_ _06867_/A vssd1 vssd1 vccd1 vccd1 _13190_/D sky130_fd_sc_hd__inv_2
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08606_ _08606_/A vssd1 vssd1 vccd1 vccd1 _08606_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_103_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09586_ _09592_/B _09583_/Y _09585_/X vssd1 vssd1 vccd1 vccd1 _09586_/Y sky130_fd_sc_hd__o21ai_1
X_06798_ _06786_/X _06790_/X _06791_/X vssd1 vssd1 vccd1 vccd1 _06798_/X sky130_fd_sc_hd__a21bo_1
XFILLER_55_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08657_/A vssd1 vssd1 vccd1 vccd1 _08642_/A sky130_fd_sc_hd__buf_2
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08468_ _13069_/Q _10390_/A _08454_/Y _12902_/Q vssd1 vssd1 vccd1 vccd1 _08468_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07419_ _11480_/X _07412_/X _13039_/Q _07415_/X vssd1 vssd1 vccd1 vccd1 _13039_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08399_ _10113_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08402_/A sky130_fd_sc_hd__or2_1
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10430_ _10433_/C vssd1 vssd1 vccd1 vccd1 _10431_/B sky130_fd_sc_hd__inv_2
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10361_ _10362_/B _10368_/D _12909_/Q _10360_/B _10350_/X vssd1 vssd1 vccd1 vccd1
+ _10361_/X sky130_fd_sc_hd__o221a_1
X_12100_ _12099_/X _12429_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _12100_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ _13081_/CLK _13080_/D _07289_/X vssd1 vssd1 vccd1 vccd1 _13080_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10292_ _10312_/A _11924_/X vssd1 vssd1 vccd1 vccd1 _10292_/Y sky130_fd_sc_hd__nor2b_4
X_12031_ _11101_/X _11099_/Y _12202_/S vssd1 vssd1 vccd1 vccd1 _12031_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12933_ _12973_/CLK _12933_/D vssd1 vssd1 vccd1 vccd1 _12933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12864_ _12864_/CLK _12864_/D _08055_/X vssd1 vssd1 vccd1 vccd1 _12864_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _11814_/X _12086_/X _11819_/S vssd1 vssd1 vccd1 vccd1 _12447_/D sky130_fd_sc_hd__mux2_1
XPHY_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _13081_/CLK _12795_/D _08379_/X vssd1 vssd1 vccd1 vccd1 _12795_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_199_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11746_ _11745_/X _11372_/X _11774_/S vssd1 vssd1 vccd1 vccd1 _12426_/D sky130_fd_sc_hd__mux2_1
XFILLER_109_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _11382_/X _09183_/A _11691_/S vssd1 vssd1 vccd1 vccd1 _11677_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10628_ _12418_/Q _12417_/Q _08926_/B vssd1 vssd1 vccd1 vccd1 _10628_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10559_ _12362_/Q vssd1 vssd1 vccd1 vccd1 _10608_/B sky130_fd_sc_hd__inv_2
XFILLER_170_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13278_ _13279_/CLK _13278_/D _06226_/X vssd1 vssd1 vccd1 vccd1 _13278_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12229_ _06283_/Y _13160_/Q _12553_/Q vssd1 vssd1 vccd1 vccd1 _12229_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07770_ _12938_/Q _11648_/S _12939_/Q _07769_/X _07569_/X vssd1 vssd1 vccd1 vccd1
+ _12939_/D sky130_fd_sc_hd__a221o_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06721_ _06719_/X _06715_/X _06720_/Y _06480_/X _13206_/Q vssd1 vssd1 vccd1 vccd1
+ _13206_/D sky130_fd_sc_hd__a32o_1
XFILLER_49_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09440_ _09440_/A vssd1 vssd1 vccd1 vccd1 _09440_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06652_ _11896_/X _06632_/B _06632_/X vssd1 vssd1 vccd1 vccd1 _06652_/X sky130_fd_sc_hd__a21bo_1
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09371_ _09359_/X _09371_/B _09371_/C _09371_/D vssd1 vssd1 vccd1 vccd1 _09371_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_75_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06583_ _06583_/A _12760_/Q vssd1 vssd1 vccd1 vccd1 _10745_/A sky130_fd_sc_hd__or2b_2
XFILLER_162_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08322_ _08325_/A vssd1 vssd1 vccd1 vccd1 _08322_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08253_ _08257_/A vssd1 vssd1 vccd1 vccd1 _08253_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_177_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07204_ _07249_/A vssd1 vssd1 vccd1 vccd1 _07204_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08184_ _08127_/Y _08128_/X _13141_/Q _10477_/A vssd1 vssd1 vccd1 vccd1 _08184_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_119_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07135_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07135_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07066_ _07078_/A vssd1 vssd1 vccd1 vccd1 _07066_/X sky130_fd_sc_hd__clkbuf_1
X_06017_ _08556_/D _06017_/B vssd1 vssd1 vccd1 vccd1 _11031_/A sky130_fd_sc_hd__or2_2
XFILLER_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07968_ _07985_/A vssd1 vssd1 vccd1 vccd1 _07968_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09707_ _13206_/Q _09706_/A _09705_/Y _09706_/Y vssd1 vssd1 vccd1 vccd1 _09708_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06919_ _06528_/X _06913_/X _06918_/Y _06841_/X _13184_/Q vssd1 vssd1 vccd1 vccd1
+ _13184_/D sky130_fd_sc_hd__a32o_1
X_07899_ _07903_/A vssd1 vssd1 vccd1 vccd1 _07899_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09638_ _09638_/A vssd1 vssd1 vccd1 vccd1 _09638_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09569_ _13155_/Q vssd1 vssd1 vccd1 vccd1 _09569_/Y sky130_fd_sc_hd__inv_2
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _10465_/X _09180_/A _11603_/S vssd1 vssd1 vccd1 vccd1 _11600_/X sky130_fd_sc_hd__mux2_1
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _12992_/CLK _12580_/D vssd1 vssd1 vccd1 vccd1 _12580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ _12820_/Q _09179_/B _11533_/S vssd1 vssd1 vccd1 vccd1 _11531_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11462_ _12905_/Q _09244_/A _11469_/S vssd1 vssd1 vccd1 vccd1 _11462_/X sky130_fd_sc_hd__mux2_1
XPHY_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13201_ _13201_/CLK _13201_/D _06767_/X vssd1 vssd1 vccd1 vccd1 _13201_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10413_ _12807_/Q _10413_/B vssd1 vssd1 vccd1 vccd1 _10415_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11393_ _09332_/A _10552_/Y _12321_/Q vssd1 vssd1 vccd1 vccd1 _11393_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13132_ _12168_/X _13132_/D _07148_/X vssd1 vssd1 vccd1 vccd1 _13132_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_3_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10344_ _10344_/A _10344_/B _10387_/A vssd1 vssd1 vccd1 vccd1 _10344_/Y sky130_fd_sc_hd__nor3_1
XFILLER_3_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13063_ _12165_/X _13063_/D _07348_/X vssd1 vssd1 vccd1 vccd1 _13063_/Q sky130_fd_sc_hd__dfrtp_1
X_10275_ _10312_/A _11923_/X vssd1 vssd1 vccd1 vccd1 _10275_/Y sky130_fd_sc_hd__nor2b_4
XFILLER_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12014_ _11118_/X _11106_/X _12201_/S vssd1 vssd1 vccd1 vccd1 _12014_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12916_ _12166_/X _12916_/D _07911_/X vssd1 vssd1 vccd1 vccd1 _12916_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12847_ _12849_/CLK _12847_/D _08098_/X vssd1 vssd1 vccd1 vccd1 _12847_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12779_/CLK _12778_/D _08425_/X vssd1 vssd1 vccd1 vccd1 _12778_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11729_ _11922_/X _11728_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _11729_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08940_ _08940_/A _08940_/B vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__nand2_4
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08871_ _08882_/A vssd1 vssd1 vccd1 vccd1 _08871_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_97_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07822_ _12893_/Q vssd1 vssd1 vccd1 vccd1 _07822_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07753_ _12940_/Q _12307_/Q _12310_/Q _07752_/Y _07616_/X vssd1 vssd1 vccd1 vccd1
+ _12940_/D sky130_fd_sc_hd__o221a_1
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06704_ _11987_/X _11990_/X _06698_/X _06699_/X _06703_/X vssd1 vssd1 vccd1 vccd1
+ _06704_/X sky130_fd_sc_hd__o32a_2
XFILLER_93_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07684_ _07684_/A _07684_/B vssd1 vssd1 vccd1 vccd1 _07685_/B sky130_fd_sc_hd__or2_1
XFILLER_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09423_ _12397_/D vssd1 vssd1 vccd1 vccd1 _09423_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06635_ _06636_/A vssd1 vssd1 vccd1 vccd1 _07019_/A sky130_fd_sc_hd__inv_2
XFILLER_52_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09354_ _12464_/Q vssd1 vssd1 vccd1 vccd1 _09354_/Y sky130_fd_sc_hd__inv_2
X_06566_ _06564_/X _06565_/X _06564_/X _06565_/X vssd1 vssd1 vccd1 vccd1 _06566_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08305_ _08128_/X _11600_/X _08307_/S vssd1 vssd1 vccd1 vccd1 _12825_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09285_ _13006_/Q _13005_/Q _09261_/X _09279_/B _09284_/X vssd1 vssd1 vccd1 vccd1
+ _09286_/B sky130_fd_sc_hd__o32a_2
XFILLER_166_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06497_ _06497_/A vssd1 vssd1 vccd1 vccd1 _06497_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08236_ _13093_/Q _10433_/A _08210_/Y _08160_/X vssd1 vssd1 vccd1 vccd1 _08237_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_166_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08167_ _12833_/Q vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__inv_2
XFILLER_147_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07118_ _07122_/A vssd1 vssd1 vccd1 vccd1 _07118_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_118_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08098_ _08098_/A vssd1 vssd1 vccd1 vccd1 _08098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07049_ _07154_/A vssd1 vssd1 vccd1 vccd1 _07063_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_122_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_148_wb_clk_i clkbuf_4_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12801_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_121_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10060_ _09484_/Y _10023_/X _10059_/Y _10025_/X vssd1 vssd1 vccd1 vccd1 _10068_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_88_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10962_ _12536_/Q vssd1 vssd1 vccd1 vccd1 _10962_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12701_ _12717_/CLK _12701_/D _08699_/X vssd1 vssd1 vccd1 vccd1 _12701_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10893_ _10864_/X _10888_/X _10836_/Y _10884_/Y _10892_/Y vssd1 vssd1 vccd1 vccd1
+ _10895_/A sky130_fd_sc_hd__o32a_2
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12632_ _13156_/CLK _12632_/D _08890_/X vssd1 vssd1 vccd1 vccd1 _12632_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ _12570_/CLK _12563_/D vssd1 vssd1 vccd1 vccd1 _12563_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11514_ _10402_/X _09184_/B _11514_/S vssd1 vssd1 vccd1 vccd1 _11514_/X sky130_fd_sc_hd__mux2_1
XPHY_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12494_ _12986_/CLK _12494_/D vssd1 vssd1 vccd1 vccd1 _12494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11445_ _12920_/Q _10794_/C _11449_/S vssd1 vssd1 vccd1 vccd1 _11445_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11376_ _11375_/X _12428_/Q _12143_/S vssd1 vssd1 vccd1 vccd1 _11376_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10327_ _07800_/X _10326_/B _10328_/B _10320_/X vssd1 vssd1 vccd1 vccd1 _10327_/X
+ sky130_fd_sc_hd__o211a_1
X_13115_ _12168_/X _13115_/D _07190_/X vssd1 vssd1 vccd1 vccd1 _13115_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13046_ _12165_/X _13046_/D _07391_/X vssd1 vssd1 vccd1 vccd1 _13046_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10258_ _10251_/Y _10038_/X _09598_/Y _10033_/X _10257_/X vssd1 vssd1 vccd1 vccd1
+ _10258_/X sky130_fd_sc_hd__o221a_2
XFILLER_140_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10189_ _10177_/Y _10134_/X _10180_/X _10188_/X vssd1 vssd1 vccd1 vccd1 _10189_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_75_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06420_ _06769_/A vssd1 vssd1 vccd1 vccd1 _06420_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06351_ _06351_/A vssd1 vssd1 vccd1 vccd1 _06351_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_175_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ _11147_/A vssd1 vssd1 vccd1 vccd1 _09070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_136_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06282_ _06075_/B _06181_/X _06075_/B _06181_/X vssd1 vssd1 vccd1 vccd1 _06283_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_147_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08021_ _08036_/A vssd1 vssd1 vccd1 vccd1 _08021_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_135_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09972_ _09972_/A vssd1 vssd1 vccd1 vccd1 _09972_/X sky130_fd_sc_hd__clkbuf_4
X_08923_ _12418_/Q vssd1 vssd1 vccd1 vccd1 _08925_/A sky130_fd_sc_hd__inv_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08854_ _08854_/A vssd1 vssd1 vccd1 vccd1 _08963_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07805_ _07801_/Y _12919_/Q _07803_/Y _07804_/X vssd1 vssd1 vccd1 vccd1 _07805_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08785_ _08784_/Y _08781_/X _06248_/X _08764_/A vssd1 vssd1 vccd1 vccd1 _12673_/D
+ sky130_fd_sc_hd__o22ai_1
X_07736_ _09475_/A vssd1 vssd1 vccd1 vccd1 _07737_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07667_ _07664_/Y _07665_/X _07666_/Y _07654_/A vssd1 vssd1 vccd1 vccd1 _07685_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09406_ _12543_/Q _10611_/B _09374_/Y _12411_/D vssd1 vssd1 vccd1 vccd1 _09406_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06618_ _12171_/X _06591_/X _12171_/X _06591_/X vssd1 vssd1 vccd1 vccd1 _06625_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_164_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07598_ _12975_/Q _12974_/Q _07598_/C vssd1 vssd1 vccd1 vccd1 _07600_/B sky130_fd_sc_hd__or3_4
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09337_ _12395_/Q vssd1 vssd1 vccd1 vccd1 _09337_/Y sky130_fd_sc_hd__inv_2
X_06549_ _06549_/A vssd1 vssd1 vccd1 vccd1 _06549_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09268_ _12299_/Q _09268_/B _09279_/D vssd1 vssd1 vccd1 vccd1 _09283_/B sky130_fd_sc_hd__and3_1
XFILLER_138_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08219_ _08193_/Y _10484_/A _08217_/Y _12826_/Q _08218_/X vssd1 vssd1 vccd1 vccd1
+ _08219_/X sky130_fd_sc_hd__o221a_1
XFILLER_194_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09199_ _09215_/A vssd1 vssd1 vccd1 vccd1 _09199_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ vssd1 vssd1 vccd1 vccd1 _11230_/HI _11230_/LO sky130_fd_sc_hd__conb_1
XFILLER_119_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11161_ vssd1 vssd1 vccd1 vccd1 _11161_/HI _11161_/LO sky130_fd_sc_hd__conb_1
XFILLER_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10112_ _12839_/Q vssd1 vssd1 vccd1 vccd1 _10112_/Y sky130_fd_sc_hd__clkinv_4
X_11092_ _10779_/X _11075_/X _06389_/X _11083_/X _11084_/X vssd1 vssd1 vccd1 vccd1
+ _11092_/X sky130_fd_sc_hd__a221o_1
XFILLER_49_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput300 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 _09071_/C sky130_fd_sc_hd__buf_1
Xinput311 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _07097_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_121_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput322 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _11966_/S sky130_fd_sc_hd__clkbuf_4
X_10043_ _10150_/A _11972_/X vssd1 vssd1 vccd1 vccd1 _10043_/Y sky130_fd_sc_hd__nor2b_1
XFILLER_76_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput333 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 input333/X sky130_fd_sc_hd__buf_2
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput344 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 _09179_/C sky130_fd_sc_hd__buf_6
XFILLER_76_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput355 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 input355/X sky130_fd_sc_hd__clkbuf_4
Xinput366 wbs_we_i vssd1 vssd1 vccd1 vccd1 _09267_/C sky130_fd_sc_hd__buf_4
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11994_ _11074_/X _11067_/X _12198_/S vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__mux2_2
XFILLER_56_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10945_ _10947_/A _10947_/B _10945_/C _10945_/D vssd1 vssd1 vccd1 vccd1 _10945_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_189_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_45_wb_clk_i clkbuf_4_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _12978_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_32_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10876_ _10876_/A vssd1 vssd1 vccd1 vccd1 _10876_/Y sky130_fd_sc_hd__inv_2
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _12942_/CLK _12616_/Q _08962_/X vssd1 vssd1 vccd1 vccd1 _12615_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12546_ _12547_/CLK _12546_/D vssd1 vssd1 vccd1 vccd1 _12546_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12477_ _12477_/CLK _12477_/D vssd1 vssd1 vccd1 vccd1 _12477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11428_ _12903_/Q _09243_/C _11433_/S vssd1 vssd1 vccd1 vccd1 _11428_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ _09329_/A _10542_/X _12321_/Q vssd1 vssd1 vccd1 vccd1 _11359_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13029_ _12164_/X _13029_/D _07441_/X vssd1 vssd1 vccd1 vccd1 _13029_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08570_ _12609_/Q _12610_/Q vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__or2_4
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07521_ _07775_/A vssd1 vssd1 vccd1 vccd1 _07522_/A sky130_fd_sc_hd__buf_2
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07452_ _07458_/A vssd1 vssd1 vccd1 vccd1 _07452_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_90_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06403_ _08504_/A vssd1 vssd1 vccd1 vccd1 _06403_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_195_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07383_ _07391_/A vssd1 vssd1 vccd1 vccd1 _07383_/X sky130_fd_sc_hd__clkbuf_1
X_09122_ _12518_/Q _09115_/X _09242_/A _09116_/X vssd1 vssd1 vccd1 vccd1 _12518_/D
+ sky130_fd_sc_hd__a22o_1
X_06334_ _06344_/A vssd1 vssd1 vccd1 vccd1 _06334_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09053_ _09058_/A _12153_/X vssd1 vssd1 vccd1 vccd1 _12564_/D sky130_fd_sc_hd__nor2b_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06265_ _06068_/X _06264_/Y _06068_/X _06264_/Y vssd1 vssd1 vccd1 vccd1 _06265_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_191_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08004_ _08004_/A vssd1 vssd1 vccd1 vccd1 _08004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_163_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06196_ _06133_/A _06070_/X _06133_/B _06070_/X _06144_/B vssd1 vssd1 vccd1 vccd1
+ _06196_/X sky130_fd_sc_hd__o221a_1
XFILLER_116_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09955_ _08767_/Y _09952_/X _06224_/X _09949_/X _09950_/X vssd1 vssd1 vccd1 vccd1
+ _09955_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_103_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08906_ _08898_/X _06332_/Y _08893_/X _12626_/Q vssd1 vssd1 vccd1 vccd1 _12626_/D
+ sky130_fd_sc_hd__o22a_1
X_09886_ _09886_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09886_/X sky130_fd_sc_hd__or2_1
XFILLER_44_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08837_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08837_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _08767_/Y _08760_/X _06224_/X _08764_/X vssd1 vssd1 vccd1 vccd1 _12678_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_72_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ _07719_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07719_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _08699_/A vssd1 vssd1 vccd1 vccd1 _08699_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ _10730_/A vssd1 vssd1 vccd1 vccd1 _10730_/X sky130_fd_sc_hd__buf_2
XPHY_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10661_ _12425_/Q vssd1 vssd1 vccd1 vccd1 _10661_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12400_ _12415_/CLK _12400_/D vssd1 vssd1 vccd1 vccd1 _12400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10592_ _10525_/A _09390_/Y _09384_/Y _10591_/Y _11403_/S vssd1 vssd1 vccd1 vccd1
+ _10592_/X sky130_fd_sc_hd__o311a_1
XFILLER_51_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12331_ _12535_/CLK _12331_/D vssd1 vssd1 vccd1 vccd1 _12331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_163_wb_clk_i clkbuf_opt_2_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _12353_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12262_ _12261_/X _12651_/Q _12618_/Q vssd1 vssd1 vccd1 vccd1 _12262_/X sky130_fd_sc_hd__mux2_2
X_11213_ vssd1 vssd1 vccd1 vccd1 _11213_/HI _11213_/LO sky130_fd_sc_hd__conb_1
XFILLER_107_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12193_ _06431_/X _11146_/A _12193_/S vssd1 vssd1 vccd1 vccd1 _12193_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11144_ _10767_/A _10737_/A _13247_/Q _10738_/A _12131_/X vssd1 vssd1 vccd1 vccd1
+ _11144_/X sky130_fd_sc_hd__a221o_1
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11075_ _11075_/A vssd1 vssd1 vccd1 vccd1 _11075_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput130 la_data_in[67] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_hd__buf_1
Xinput141 la_data_in[77] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_hd__buf_1
Xinput152 la_data_in[87] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_hd__buf_1
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10026_ _10022_/Y _10023_/X _10024_/Y _10025_/X vssd1 vssd1 vccd1 vccd1 _10041_/B
+ sky130_fd_sc_hd__o22a_1
Xinput163 la_data_in[97] vssd1 vssd1 vccd1 vccd1 input163/X sky130_fd_sc_hd__buf_1
XFILLER_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput174 la_oenb[106] vssd1 vssd1 vccd1 vccd1 input174/X sky130_fd_sc_hd__buf_1
XFILLER_110_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput185 la_oenb[116] vssd1 vssd1 vccd1 vccd1 input185/X sky130_fd_sc_hd__buf_1
Xinput196 la_oenb[126] vssd1 vssd1 vccd1 vccd1 input196/X sky130_fd_sc_hd__buf_1
XFILLER_64_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11977_ _10149_/Y _12793_/Q _11981_/S vssd1 vssd1 vccd1 vccd1 _11977_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10928_ _12531_/Q vssd1 vssd1 vccd1 vccd1 _10930_/A sky130_fd_sc_hd__inv_2
XFILLER_177_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10859_ _10859_/A vssd1 vssd1 vccd1 vccd1 _10859_/Y sky130_fd_sc_hd__inv_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12529_ _12529_/CLK _12529_/D vssd1 vssd1 vccd1 vccd1 _12529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06050_ _12740_/Q _12708_/Q _12740_/Q _12708_/Q vssd1 vssd1 vccd1 vccd1 _06050_/X
+ sky130_fd_sc_hd__o2bb2a_1
Xoutput604 _12290_/Q vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09740_ _09740_/A vssd1 vssd1 vccd1 vccd1 _09740_/Y sky130_fd_sc_hd__inv_2
X_06952_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06952_/X sky130_fd_sc_hd__clkbuf_1
.ends

